module IOB(
  input  [31:0] io_in_0,
  output [31:0] io_out_0
);
  assign io_out_0 = io_in_0; // @[IOB.scala 66:42]
endmodule
module Muxn(
  input         io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out
);
  assign io_out = io_config ? io_in_1 : io_in_0; // @[Multiplexer.scala 20:10]
endmodule
module ConfigMem(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output        io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  configmem_0_0; // @[ConfigMem.scala 81:26]
  wire  _GEN_0 = io_cfg_en & io_cfg_data[0]; // @[ConfigMem.scala 111:54]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  configmem_0_0 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 1'h0;
    end else if (io_cfg_en) begin
      configmem_0_0 <= _GEN_0;
    end
  end
endmodule
module IOB_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'h6 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module IOB_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'h7 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module IOB_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'h8 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module IOB_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'hd3 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module IOB_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'hd4 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module IOB_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_0; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_in_1; // @[IOB.scala 46:41]
  wire [31:0] Muxn_io_out; // @[IOB.scala 46:41]
  wire  ConfigMem_clock; // @[IOB.scala 47:21]
  wire  ConfigMem_reset; // @[IOB.scala 47:21]
  wire  ConfigMem_io_cfg_en; // @[IOB.scala 47:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[IOB.scala 47:21]
  wire  ConfigMem_io_out_0; // @[IOB.scala 47:21]
  wire  _T_1 = 10'hd5 == io_cfg_addr[13:4]; // @[IOB.scala 48:50]
  Muxn Muxn ( // @[IOB.scala 46:41]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  ConfigMem ConfigMem ( // @[IOB.scala 47:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  assign io_out_0 = Muxn_io_out; // @[IOB.scala 61:17]
  assign Muxn_io_config = ConfigMem_io_out_0; // @[IOB.scala 62:22]
  assign Muxn_io_in_0 = io_in_0; // @[IOB.scala 59:23]
  assign Muxn_io_in_1 = io_in_1; // @[IOB.scala 59:23]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[IOB.scala 48:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[IOB.scala 53:21]
endmodule
module ALU(
  input  [4:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out
);
  wire [31:0] _T_4 = io_in_0 + io_in_1; // @[Operations.scala 131:41]
  wire [31:0] _T_8 = io_in_0 - io_in_1; // @[Operations.scala 133:41]
  wire [63:0] _T_11 = io_in_0 * io_in_1; // @[Operations.scala 135:41]
  wire [31:0] _T_14 = io_in_0 & io_in_1; // @[Operations.scala 146:41]
  wire [31:0] _T_17 = io_in_0 | io_in_1; // @[Operations.scala 148:41]
  wire [31:0] _T_20 = io_in_0 ^ io_in_1; // @[Operations.scala 150:41]
  wire  _T_21 = 5'h0 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_22 = _T_21 ? io_in_0 : 32'h0; // @[Mux.scala 80:57]
  wire  _T_23 = 5'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_24 = _T_23 ? _T_4 : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 5'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_26 = _T_25 ? _T_8 : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 5'h3 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_28 = _T_27 ? _T_11 : {{32'd0}, _T_26}; // @[Mux.scala 80:57]
  wire  _T_29 = 5'h4 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_30 = _T_29 ? {{32'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 5'h5 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_32 = _T_31 ? {{32'd0}, _T_17} : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 5'h6 == io_config; // @[Mux.scala 80:60]
  wire [63:0] _T_34 = _T_33 ? {{32'd0}, _T_20} : _T_32; // @[Mux.scala 80:57]
  assign io_out = _T_34[31:0]; // @[ALU.scala 25:10]
endmodule
module RF(
  input         clock,
  input         reset,
  input         io_en,
  input  [31:0] io_in_0,
  output [31:0] io_out_0,
  output [31:0] io_out_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[RegFile.scala 24:21]
  assign io_out_0 = regs_0; // @[RegFile.scala 37:42]
  assign io_out_1 = regs_0; // @[RegFile.scala 37:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (io_en) begin
      regs_0 <= io_in_0;
    end
  end
endmodule
module DelayPipe(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_config,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[DelayPipe.scala 70:21]
  reg [31:0] regs_1; // @[DelayPipe.scala 70:21]
  reg [31:0] regs_2; // @[DelayPipe.scala 70:21]
  reg [31:0] regs_3; // @[DelayPipe.scala 70:21]
  reg [31:0] regs_4; // @[DelayPipe.scala 70:21]
  reg [2:0] wptr; // @[DelayPipe.scala 71:21]
  reg [2:0] rptr; // @[DelayPipe.scala 72:21]
  reg [2:0] config_temp; // @[DelayPipe.scala 74:28]
  wire  _T_1 = wptr < 3'h4; // @[DelayPipe.scala 77:23]
  wire  _T_2 = io_en & _T_1; // @[DelayPipe.scala 77:14]
  wire [2:0] _T_4 = wptr + 3'h1; // @[DelayPipe.scala 78:17]
  wire  _T_7 = _T_4 >= io_config; // @[DelayPipe.scala 83:17]
  wire [2:0] _T_11 = _T_4 - io_config; // @[DelayPipe.scala 84:24]
  wire [2:0] _T_13 = 3'h6 + wptr; // @[DelayPipe.scala 86:30]
  wire [2:0] _T_15 = _T_13 - io_config; // @[DelayPipe.scala 86:37]
  wire  _T_16 = io_config > 3'h0; // @[DelayPipe.scala 90:28]
  wire  _T_17 = io_en & _T_16; // @[DelayPipe.scala 90:14]
  reg [2:0] cnt; // @[DelayPipe.scala 94:20]
  wire  _T_18 = ~io_en; // @[DelayPipe.scala 95:8]
  wire  _T_19 = config_temp != io_config; // @[DelayPipe.scala 97:26]
  wire  _T_20 = cnt < io_config; // @[DelayPipe.scala 99:18]
  wire [2:0] _T_22 = cnt + 3'h1; // @[DelayPipe.scala 100:16]
  wire  _T_23 = 3'h0 == io_config; // @[DelayPipe.scala 103:22]
  wire  _T_24 = io_en & _T_23; // @[DelayPipe.scala 103:14]
  wire  _T_25 = cnt == io_config; // @[DelayPipe.scala 105:28]
  wire  _T_26 = io_en & _T_25; // @[DelayPipe.scala 105:20]
  wire [31:0] _GEN_16 = 3'h1 == rptr ? regs_1 : regs_0; // @[DelayPipe.scala 106:12]
  wire [31:0] _GEN_17 = 3'h2 == rptr ? regs_2 : _GEN_16; // @[DelayPipe.scala 106:12]
  wire [31:0] _GEN_18 = 3'h3 == rptr ? regs_3 : _GEN_17; // @[DelayPipe.scala 106:12]
  wire [31:0] _GEN_19 = 3'h4 == rptr ? regs_4 : _GEN_18; // @[DelayPipe.scala 106:12]
  wire [31:0] _GEN_20 = _T_26 ? _GEN_19 : 32'h0; // @[DelayPipe.scala 105:43]
  assign io_out = _T_24 ? io_in : _GEN_20; // @[DelayPipe.scala 104:12 DelayPipe.scala 106:12 DelayPipe.scala 108:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  wptr = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  rptr = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  config_temp = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  cnt = _RAND_8[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (_T_17) begin
      if (3'h0 == wptr) begin
        regs_0 <= io_in;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else if (_T_17) begin
      if (3'h1 == wptr) begin
        regs_1 <= io_in;
      end
    end
    if (reset) begin
      regs_2 <= 32'h0;
    end else if (_T_17) begin
      if (3'h2 == wptr) begin
        regs_2 <= io_in;
      end
    end
    if (reset) begin
      regs_3 <= 32'h0;
    end else if (_T_17) begin
      if (3'h3 == wptr) begin
        regs_3 <= io_in;
      end
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else if (_T_17) begin
      if (3'h4 == wptr) begin
        regs_4 <= io_in;
      end
    end
    if (reset) begin
      wptr <= 3'h0;
    end else if (_T_2) begin
      wptr <= _T_4;
    end else begin
      wptr <= 3'h0;
    end
    if (reset) begin
      rptr <= 3'h0;
    end else if (_T_7) begin
      rptr <= _T_11;
    end else begin
      rptr <= _T_15;
    end
    if (reset) begin
      config_temp <= 3'h0;
    end else begin
      config_temp <= io_config;
    end
    if (reset) begin
      cnt <= 3'h0;
    end else if (_T_18) begin
      cnt <= 3'h0;
    end else if (_T_19) begin
      cnt <= 3'h1;
    end else if (_T_20) begin
      cnt <= _T_22;
    end
  end
endmodule
module Muxn_6(
  input  [2:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  output [31:0] io_out
);
  wire  _T_2 = 3'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 3'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_5 = _T_4 ? io_in_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 3'h3 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_7 = _T_6 ? io_in_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 3'h4 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_9 = _T_8 ? io_in_4 : _T_7; // @[Mux.scala 80:57]
  wire  _T_10 = 3'h5 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_10 ? io_in_5 : _T_9; // @[Multiplexer.scala 20:10]
endmodule
module ConfigMem_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input         io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [48:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [48:0] configmem_0_0; // @[ConfigMem.scala 81:26]
  wire  _T_1 = ~io_cfg_addr; // @[ConfigMem.scala 120:38]
  wire  _T_2 = io_cfg_en & _T_1; // @[ConfigMem.scala 120:22]
  wire [48:0] _T_4 = {configmem_0_0[48:32],io_cfg_data}; // @[Cat.scala 29:58]
  wire [48:0] _GEN_0 = _T_2 ? _T_4 : configmem_0_0; // @[ConfigMem.scala 120:47]
  wire  _T_6 = io_cfg_en & io_cfg_addr; // @[ConfigMem.scala 120:22]
  wire [63:0] _T_8 = {io_cfg_data,configmem_0_0[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_1 = _T_6 ? _T_8 : {{15'd0}, _GEN_0}; // @[ConfigMem.scala 120:47]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  configmem_0_0 = _RAND_0[48:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 49'h0;
    end else begin
      configmem_0_0 <= _GEN_1[48:0];
    end
  end
endmodule
module GPE(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h11 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_1(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h12 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_2(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h13 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_3(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h1b == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_4(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h1c == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_5(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h1d == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h25 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h26 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h27 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h2f == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h30 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h31 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_12(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h39 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_13(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h3a == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_14(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h3b == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_15(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h43 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h44 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h45 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h4d == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h4e == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h4f == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h57 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h58 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h59 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h61 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h62 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h63 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h6b == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h6c == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h6d == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h75 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h76 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_32(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h77 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_33(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h7f == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_34(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h80 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_35(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h81 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_36(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h89 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_37(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h8a == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_38(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h8b == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_39(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h93 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_40(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h94 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_41(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h95 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_42(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h9d == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_43(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h9e == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_44(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'h9f == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_45(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'ha7 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_46(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'ha8 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_47(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'ha9 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_48(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hb1 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_49(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hb2 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_50(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hb3 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_51(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hbb == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_52(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hbc == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_53(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hbd == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_54(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hc5 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_55(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hc6 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module GPE_56(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  input  [31:0] io_in_6,
  input  [31:0] io_in_7,
  output [31:0] io_out_0
);
  wire [4:0] alu_io_config; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_0; // @[PE.scala 52:19]
  wire [31:0] alu_io_in_1; // @[PE.scala 52:19]
  wire [31:0] alu_io_out; // @[PE.scala 52:19]
  wire  rf_clock; // @[PE.scala 53:18]
  wire  rf_reset; // @[PE.scala 53:18]
  wire  rf_io_en; // @[PE.scala 53:18]
  wire [31:0] rf_io_in_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_0; // @[PE.scala 53:18]
  wire [31:0] rf_io_out_1; // @[PE.scala 53:18]
  wire  DelayPipe_clock; // @[PE.scala 54:54]
  wire  DelayPipe_reset; // @[PE.scala 54:54]
  wire  DelayPipe_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_io_out; // @[PE.scala 54:54]
  wire  DelayPipe_1_clock; // @[PE.scala 54:54]
  wire  DelayPipe_1_reset; // @[PE.scala 54:54]
  wire  DelayPipe_1_io_en; // @[PE.scala 54:54]
  wire [2:0] DelayPipe_1_io_config; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_in; // @[PE.scala 54:54]
  wire [31:0] DelayPipe_1_io_out; // @[PE.scala 54:54]
  wire [2:0] Muxn_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_io_out; // @[PE.scala 57:49]
  wire [2:0] Muxn_1_io_config; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_0; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_1; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_2; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_3; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_4; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_in_5; // @[PE.scala 57:49]
  wire [31:0] Muxn_1_io_out; // @[PE.scala 57:49]
  wire  cfg_clock; // @[PE.scala 98:19]
  wire  cfg_reset; // @[PE.scala 98:19]
  wire  cfg_io_cfg_en; // @[PE.scala 98:19]
  wire  cfg_io_cfg_addr; // @[PE.scala 98:19]
  wire [31:0] cfg_io_cfg_data; // @[PE.scala 98:19]
  wire [48:0] cfg_io_out_0; // @[PE.scala 98:19]
  wire  _T_1 = 10'hc7 == io_cfg_addr[13:4]; // @[PE.scala 99:48]
  wire [48:0] cfgOut = cfg_io_out_0; // @[PE.scala 108:20 PE.scala 109:10]
  ALU alu ( // @[PE.scala 52:19]
    .io_config(alu_io_config),
    .io_in_0(alu_io_in_0),
    .io_in_1(alu_io_in_1),
    .io_out(alu_io_out)
  );
  RF rf ( // @[PE.scala 53:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_en(rf_io_en),
    .io_in_0(rf_io_in_0),
    .io_out_0(rf_io_out_0),
    .io_out_1(rf_io_out_1)
  );
  DelayPipe DelayPipe ( // @[PE.scala 54:54]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[PE.scala 54:54]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  Muxn_6 Muxn ( // @[PE.scala 57:49]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_in_4(Muxn_io_in_4),
    .io_in_5(Muxn_io_in_5),
    .io_out(Muxn_io_out)
  );
  Muxn_6 Muxn_1 ( // @[PE.scala 57:49]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_in_4(Muxn_1_io_in_4),
    .io_in_5(Muxn_1_io_in_5),
    .io_out(Muxn_1_io_out)
  );
  ConfigMem_6 cfg ( // @[PE.scala 98:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_out_0 = rf_io_out_0; // @[PE.scala 79:13]
  assign alu_io_config = cfgOut[36:32]; // @[PE.scala 112:19]
  assign alu_io_in_0 = DelayPipe_io_out; // @[PE.scala 73:18]
  assign alu_io_in_1 = DelayPipe_1_io_out; // @[PE.scala 73:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_en = io_en; // @[PE.scala 77:12]
  assign rf_io_in_0 = alu_io_out; // @[PE.scala 78:15]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_io_config = cfgOut[39:37]; // @[PE.scala 125:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[PE.scala 72:23]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[PE.scala 71:23]
  assign DelayPipe_1_io_config = cfgOut[42:40]; // @[PE.scala 125:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[PE.scala 72:23]
  assign Muxn_io_config = cfgOut[45:43]; // @[PE.scala 133:23]
  assign Muxn_io_in_0 = io_in_0; // @[PE.scala 64:12]
  assign Muxn_io_in_1 = io_in_1; // @[PE.scala 64:12]
  assign Muxn_io_in_2 = io_in_2; // @[PE.scala 64:12]
  assign Muxn_io_in_3 = io_in_3; // @[PE.scala 64:12]
  assign Muxn_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign Muxn_1_io_config = cfgOut[48:46]; // @[PE.scala 133:23]
  assign Muxn_1_io_in_0 = io_in_4; // @[PE.scala 64:12]
  assign Muxn_1_io_in_1 = io_in_5; // @[PE.scala 64:12]
  assign Muxn_1_io_in_2 = io_in_6; // @[PE.scala 64:12]
  assign Muxn_1_io_in_3 = io_in_7; // @[PE.scala 64:12]
  assign Muxn_1_io_in_4 = cfgOut[31:0]; // @[PE.scala 66:12]
  assign Muxn_1_io_in_5 = rf_io_out_1; // @[PE.scala 68:12]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_1; // @[PE.scala 99:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[PE.scala 100:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[PE.scala 104:19]
endmodule
module ConfigMem_63(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [17:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] configmem_0_0; // @[ConfigMem.scala 81:26]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  configmem_0_0 = _RAND_0[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 18'h0;
    end else if (io_cfg_en) begin
      if (io_cfg_en) begin
        configmem_0_0 <= io_cfg_data[17:0];
      end else begin
        configmem_0_0 <= 18'h0;
      end
    end
  end
endmodule
module Muxn_120(
  input  [1:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  output [31:0] io_out
);
  wire  _T_2 = 2'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h2 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_4 ? io_in_2 : _T_3; // @[Multiplexer.scala 20:10]
endmodule
module Muxn_124(
  input  [2:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  output [31:0] io_out
);
  wire  _T_2 = 3'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_4 = 3'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_5 = _T_4 ? io_in_2 : _T_3; // @[Mux.scala 80:57]
  wire  _T_6 = 3'h3 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_7 = _T_6 ? io_in_3 : _T_5; // @[Mux.scala 80:57]
  wire  _T_8 = 3'h4 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_8 ? io_in_4 : _T_7; // @[Multiplexer.scala 20:10]
endmodule
module Muxn_126(
  input  [1:0]  io_config,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  output [31:0] io_out
);
  wire  _T = 2'h1 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? io_in_1 : io_in_0; // @[Mux.scala 80:57]
  wire  _T_2 = 2'h2 == io_config; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? io_in_2 : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h3 == io_config; // @[Mux.scala 80:60]
  assign io_out = _T_4 ? io_in_3 : _T_3; // @[Multiplexer.scala 20:10]
endmodule
module GIB(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [17:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hb == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_63 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_124 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_124 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_in_4(Muxn_5_io_in_4),
    .io_out(Muxn_5_io_out)
  );
  Muxn_126 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_126 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNE_0 = Muxn_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_1_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_2_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_3_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_6_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_7_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[10:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[13:11]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:16]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module ConfigMem_64(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [23:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] configmem_0_0; // @[ConfigMem.scala 81:26]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  configmem_0_0 = _RAND_0[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 24'h0;
    end else if (io_cfg_en) begin
      if (io_cfg_en) begin
        configmem_0_0 <= io_cfg_data[23:0];
      end else begin
        configmem_0_0 <= 24'h0;
      end
    end
  end
endmodule
module GIB_1(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hc == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_126 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_2(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hd == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_126 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_in_3(Muxn_1_io_in_3),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_2_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_3(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [17:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'he == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_10; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  ConfigMem_63 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_126 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_124 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_in_4(Muxn_5_io_in_4),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_126 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_1_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_2_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_3_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_10; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_16; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[12:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[15:13]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:16]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_10 <= Muxn_4_io_out;
    _T_16 <= Muxn_7_io_out;
  end
endmodule
module GIB_4(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h15 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module ConfigMem_68(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [31:0] io_cfg_data,
  output [27:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [27:0] configmem_0_0; // @[ConfigMem.scala 81:26]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  configmem_0_0 = _RAND_0[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 28'h0;
    end else if (io_cfg_en) begin
      if (io_cfg_en) begin
        configmem_0_0 <= io_cfg_data[27:0];
      end else begin
        configmem_0_0 <= 28'h0;
      end
    end
  end
endmodule
module GIB_5(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h16 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h17 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h18 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h1f == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h20 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h21 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h22 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_12(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h29 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_13(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h2a == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_14(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h2b == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_15(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h2c == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h33 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h34 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h35 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h36 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h3d == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h3e == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h3f == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h40 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h47 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h48 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h49 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h4a == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h51 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h52 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h53 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h54 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_32(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h5b == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_33(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h5c == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_34(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h5d == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_35(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h5e == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_36(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h65 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_37(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h66 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_38(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h67 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_39(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h68 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_40(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h6f == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_41(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h70 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_42(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h71 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_43(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h72 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_44(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h79 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_45(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h7a == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_46(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h7b == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_47(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h7c == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_48(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h83 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_49(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h84 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_50(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h85 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_51(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h86 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_52(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h8d == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_53(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h8e == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_54(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h8f == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_55(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h90 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_56(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h97 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_57(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h98 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_58(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h99 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_59(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'h9a == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_60(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'ha1 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_61(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'ha2 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_62(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'ha3 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_63(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'ha4 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_64(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hab == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_65(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hac == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_66(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'had == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_67(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hae == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_68(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hb5 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_69(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hb6 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_70(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hb7 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_71(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hb8 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module GIB_72(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hbf == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_126 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_in_3(Muxn_io_in_3),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_9_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_73(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hc0 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  reg [31:0] _T_20; // @[Interconnect.scala 617:55]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_14; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_16; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_18; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_20; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_14 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_16 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_14 <= Muxn_8_io_out;
    _T_16 <= Muxn_9_io_out;
    _T_18 <= Muxn_10_io_out;
    _T_20 <= Muxn_11_io_out;
  end
endmodule
module GIB_74(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  output [31:0] io_ipinSE_1,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [27:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_10_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_10_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_11_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_11_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hc1 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_68 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_120 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_out(Muxn_6_io_out)
  );
  Muxn_120 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  Muxn_124 Muxn_10 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_10_io_config),
    .io_in_0(Muxn_10_io_in_0),
    .io_in_1(Muxn_10_io_in_1),
    .io_in_2(Muxn_10_io_in_2),
    .io_in_3(Muxn_10_io_in_3),
    .io_in_4(Muxn_10_io_in_4),
    .io_out(Muxn_10_io_out)
  );
  Muxn_124 Muxn_11 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_11_io_config),
    .io_in_0(Muxn_11_io_in_0),
    .io_in_1(Muxn_11_io_in_1),
    .io_in_2(Muxn_11_io_in_2),
    .io_in_3(Muxn_11_io_in_3),
    .io_in_4(Muxn_11_io_in_4),
    .io_out(Muxn_11_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSE_1 = Muxn_5_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_6_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_7_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_8_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_9_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_10_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign io_otrackS_0 = Muxn_11_io_out; // @[Interconnect.scala 564:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[13:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[15:14]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[18:16]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[21:19]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_config = ConfigMem_io_out_0[24:22]; // @[Interconnect.scala 623:23]
  assign Muxn_10_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_10_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_config = ConfigMem_io_out_0[27:25]; // @[Interconnect.scala 623:23]
  assign Muxn_11_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_11_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_75(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  output [31:0] io_ipinSW_1,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackS_0,
  output [31:0] io_otrackS_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hc2 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_18; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_126 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_in_3(Muxn_2_io_in_3),
    .io_out(Muxn_2_io_out)
  );
  Muxn_126 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_in_3(Muxn_3_io_in_3),
    .io_out(Muxn_3_io_out)
  );
  Muxn_120 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_out(Muxn_4_io_out)
  );
  Muxn_120 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_4_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_ipinSW_1 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackS_0 = _T_18; // @[Interconnect.scala 564:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_3 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = io_itrackS_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_18 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_18 <= Muxn_9_io_out;
  end
endmodule
module GIB_76(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [17:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hc9 == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  ConfigMem_63 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_124 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_in_4(Muxn_4_io_in_4),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_126 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_1_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_3_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_otrackN_0 = _T_12; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_14; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[10:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[12:11]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:13]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_5_io_out;
    _T_14 <= Muxn_6_io_out;
  end
endmodule
module GIB_77(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hca == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_126 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_6_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_7_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign io_otrackE_0 = Muxn_8_io_out; // @[Interconnect.scala 563:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
endmodule
module GIB_78(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  output [31:0] io_ipinNE_1,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSE_0,
  input  [31:0] io_opinSE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0,
  input  [31:0] io_itrackE_0,
  output [31:0] io_otrackE_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [23:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_8_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_8_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_9_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_9_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hcb == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  reg [31:0] _T_12; // @[Interconnect.scala 617:55]
  reg [31:0] _T_14; // @[Interconnect.scala 617:55]
  reg [31:0] _T_16; // @[Interconnect.scala 617:55]
  ConfigMem_64 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_126 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  Muxn_124 Muxn_8 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_8_io_config),
    .io_in_0(Muxn_8_io_in_0),
    .io_in_1(Muxn_8_io_in_1),
    .io_in_2(Muxn_8_io_in_2),
    .io_in_3(Muxn_8_io_in_3),
    .io_in_4(Muxn_8_io_in_4),
    .io_out(Muxn_8_io_out)
  );
  Muxn_124 Muxn_9 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_9_io_config),
    .io_in_0(Muxn_9_io_in_0),
    .io_in_1(Muxn_9_io_in_1),
    .io_in_2(Muxn_9_io_in_2),
    .io_in_3(Muxn_9_io_in_3),
    .io_in_4(Muxn_9_io_in_4),
    .io_out(Muxn_9_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinNE_1 = Muxn_3_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSE_0 = Muxn_4_io_out; // @[Interconnect.scala 560:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_5_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = _T_12; // @[Interconnect.scala 561:21 Interconnect.scala 617:45]
  assign io_otrackN_0 = _T_14; // @[Interconnect.scala 562:21 Interconnect.scala 617:45]
  assign io_otrackE_0 = _T_16; // @[Interconnect.scala 563:21 Interconnect.scala 617:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinSE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_config = ConfigMem_io_out_0[20:18]; // @[Interconnect.scala 623:23]
  assign Muxn_8_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_8_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_config = ConfigMem_io_out_0[23:21]; // @[Interconnect.scala 623:23]
  assign Muxn_9_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_9_io_in_4 = io_itrackE_0; // @[Interconnect.scala 615:63]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_16 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_12 <= Muxn_6_io_out;
    _T_14 <= Muxn_7_io_out;
    _T_16 <= Muxn_8_io_out;
  end
endmodule
module GIB_79(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [31:0] io_ipinNW_0,
  output [31:0] io_ipinNW_1,
  input  [31:0] io_opinNW_0,
  output [31:0] io_ipinNE_0,
  input  [31:0] io_opinNE_0,
  output [31:0] io_ipinSW_0,
  input  [31:0] io_opinSW_0,
  input  [31:0] io_itrackW_0,
  output [31:0] io_otrackW_0,
  input  [31:0] io_itrackN_0,
  output [31:0] io_otrackN_0
);
  wire  ConfigMem_clock; // @[Interconnect.scala 601:21]
  wire  ConfigMem_reset; // @[Interconnect.scala 601:21]
  wire  ConfigMem_io_cfg_en; // @[Interconnect.scala 601:21]
  wire [31:0] ConfigMem_io_cfg_data; // @[Interconnect.scala 601:21]
  wire [17:0] ConfigMem_io_out_0; // @[Interconnect.scala 601:21]
  wire [1:0] Muxn_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_1_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_1_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_2_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_2_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_3_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_3_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_4_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_4_io_out; // @[Interconnect.scala 613:25]
  wire [1:0] Muxn_5_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_5_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_6_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_6_io_out; // @[Interconnect.scala 613:25]
  wire [2:0] Muxn_7_io_config; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_0; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_1; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_2; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_3; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_in_4; // @[Interconnect.scala 613:25]
  wire [31:0] Muxn_7_io_out; // @[Interconnect.scala 613:25]
  wire  _T_1 = 10'hcc == io_cfg_addr[13:4]; // @[Interconnect.scala 602:50]
  ConfigMem_63 ConfigMem ( // @[Interconnect.scala 601:21]
    .clock(ConfigMem_clock),
    .reset(ConfigMem_reset),
    .io_cfg_en(ConfigMem_io_cfg_en),
    .io_cfg_data(ConfigMem_io_cfg_data),
    .io_out_0(ConfigMem_io_out_0)
  );
  Muxn_120 Muxn ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_in_2(Muxn_io_in_2),
    .io_out(Muxn_io_out)
  );
  Muxn_120 Muxn_1 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_in_2(Muxn_1_io_in_2),
    .io_out(Muxn_1_io_out)
  );
  Muxn_120 Muxn_2 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_2_io_config),
    .io_in_0(Muxn_2_io_in_0),
    .io_in_1(Muxn_2_io_in_1),
    .io_in_2(Muxn_2_io_in_2),
    .io_out(Muxn_2_io_out)
  );
  Muxn_120 Muxn_3 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_3_io_config),
    .io_in_0(Muxn_3_io_in_0),
    .io_in_1(Muxn_3_io_in_1),
    .io_in_2(Muxn_3_io_in_2),
    .io_out(Muxn_3_io_out)
  );
  Muxn_126 Muxn_4 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_4_io_config),
    .io_in_0(Muxn_4_io_in_0),
    .io_in_1(Muxn_4_io_in_1),
    .io_in_2(Muxn_4_io_in_2),
    .io_in_3(Muxn_4_io_in_3),
    .io_out(Muxn_4_io_out)
  );
  Muxn_126 Muxn_5 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_5_io_config),
    .io_in_0(Muxn_5_io_in_0),
    .io_in_1(Muxn_5_io_in_1),
    .io_in_2(Muxn_5_io_in_2),
    .io_in_3(Muxn_5_io_in_3),
    .io_out(Muxn_5_io_out)
  );
  Muxn_124 Muxn_6 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_6_io_config),
    .io_in_0(Muxn_6_io_in_0),
    .io_in_1(Muxn_6_io_in_1),
    .io_in_2(Muxn_6_io_in_2),
    .io_in_3(Muxn_6_io_in_3),
    .io_in_4(Muxn_6_io_in_4),
    .io_out(Muxn_6_io_out)
  );
  Muxn_124 Muxn_7 ( // @[Interconnect.scala 613:25]
    .io_config(Muxn_7_io_config),
    .io_in_0(Muxn_7_io_in_0),
    .io_in_1(Muxn_7_io_in_1),
    .io_in_2(Muxn_7_io_in_2),
    .io_in_3(Muxn_7_io_in_3),
    .io_in_4(Muxn_7_io_in_4),
    .io_out(Muxn_7_io_out)
  );
  assign io_ipinNW_0 = Muxn_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNW_1 = Muxn_1_io_out; // @[Interconnect.scala 557:20 Interconnect.scala 619:45]
  assign io_ipinNE_0 = Muxn_2_io_out; // @[Interconnect.scala 558:20 Interconnect.scala 619:45]
  assign io_ipinSW_0 = Muxn_3_io_out; // @[Interconnect.scala 559:20 Interconnect.scala 619:45]
  assign io_otrackW_0 = Muxn_4_io_out; // @[Interconnect.scala 561:21 Interconnect.scala 619:45]
  assign io_otrackN_0 = Muxn_5_io_out; // @[Interconnect.scala 562:21 Interconnect.scala 619:45]
  assign ConfigMem_clock = clock;
  assign ConfigMem_reset = reset;
  assign ConfigMem_io_cfg_en = io_cfg_en & _T_1; // @[Interconnect.scala 602:19]
  assign ConfigMem_io_cfg_data = io_cfg_data; // @[Interconnect.scala 607:21]
  assign Muxn_io_config = ConfigMem_io_out_0[1:0]; // @[Interconnect.scala 623:23]
  assign Muxn_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_config = ConfigMem_io_out_0[3:2]; // @[Interconnect.scala 623:23]
  assign Muxn_1_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_1 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_1_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_config = ConfigMem_io_out_0[5:4]; // @[Interconnect.scala 623:23]
  assign Muxn_2_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_2_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_config = ConfigMem_io_out_0[7:6]; // @[Interconnect.scala 623:23]
  assign Muxn_3_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_3_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_config = ConfigMem_io_out_0[9:8]; // @[Interconnect.scala 623:23]
  assign Muxn_4_io_in_0 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_1 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_4_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_config = ConfigMem_io_out_0[11:10]; // @[Interconnect.scala 623:23]
  assign Muxn_5_io_in_0 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_1 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_2 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_5_io_in_3 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_config = ConfigMem_io_out_0[14:12]; // @[Interconnect.scala 623:23]
  assign Muxn_6_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_1 = io_opinSW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_6_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_config = ConfigMem_io_out_0[17:15]; // @[Interconnect.scala 623:23]
  assign Muxn_7_io_in_0 = io_opinNW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_1 = io_opinNE_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_2 = io_itrackW_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_3 = io_itrackN_0; // @[Interconnect.scala 615:63]
  assign Muxn_7_io_in_4 = 32'h0; // @[Interconnect.scala 615:63]
endmodule
module single_port_ram(
  input         clock,
  input         io_enable,
  input         io_write_enable,
  input  [5:0]  io_addr,
  input  [31:0] io_dataIn,
  output [31:0] io_dataOut
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:63]; // @[SRAM.scala 125:24]
  wire [31:0] mem__T_r_data; // @[SRAM.scala 125:24]
  wire [5:0] mem__T_r_addr; // @[SRAM.scala 125:24]
  wire [31:0] mem__T_w_data; // @[SRAM.scala 125:24]
  wire [5:0] mem__T_w_addr; // @[SRAM.scala 125:24]
  wire  mem__T_w_mask; // @[SRAM.scala 125:24]
  wire  mem__T_w_en; // @[SRAM.scala 125:24]
  reg  mem__T_r_en_pipe_0;
  reg [5:0] mem__T_r_addr_pipe_0;
  wire  _GEN_8 = io_enable & io_write_enable; // @[SRAM.scala 127:19]
  wire  _GEN_11 = ~_GEN_8;
  assign mem__T_r_addr = mem__T_r_addr_pipe_0;
  assign mem__T_r_data = mem[mem__T_r_addr]; // @[SRAM.scala 125:24]
  assign mem__T_w_data = io_dataIn;
  assign mem__T_w_addr = io_addr;
  assign mem__T_w_mask = io_write_enable;
  assign mem__T_w_en = io_enable & _GEN_8;
  assign io_dataOut = mem__T_r_data; // @[SRAM.scala 130:34]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem__T_r_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_w_en & mem__T_w_mask) begin
      mem[mem__T_w_addr] <= mem__T_w_data; // @[SRAM.scala 125:24]
    end
    mem__T_r_en_pipe_0 <= io_enable & _GEN_11;
    if (io_enable & _GEN_11) begin
      mem__T_r_addr_pipe_0 <= io_addr;
    end
  end
endmodule
module ConfigMem_143(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input         io_cfg_addr,
  input  [31:0] io_cfg_data,
  output [40:0] io_out_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [40:0] configmem_0_0; // @[ConfigMem.scala 81:26]
  wire  _T_1 = ~io_cfg_addr; // @[ConfigMem.scala 120:38]
  wire  _T_2 = io_cfg_en & _T_1; // @[ConfigMem.scala 120:22]
  wire [40:0] _T_4 = {configmem_0_0[40:32],io_cfg_data}; // @[Cat.scala 29:58]
  wire [40:0] _GEN_0 = _T_2 ? _T_4 : configmem_0_0; // @[ConfigMem.scala 120:47]
  wire  _T_6 = io_cfg_en & io_cfg_addr; // @[ConfigMem.scala 120:22]
  wire [63:0] _T_8 = {io_cfg_data,configmem_0_0[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_1 = _T_6 ? _T_8 : {{23'd0}, _GEN_0}; // @[ConfigMem.scala 120:47]
  assign io_out_0 = configmem_0_0; // @[ConfigMem.scala 140:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  configmem_0_0 = _RAND_0[40:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      configmem_0_0 <= 41'h0;
    end else begin
      configmem_0_0 <= _GEN_1[40:0];
    end
  end
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h10 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_1(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h14 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_2(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h1a == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_3(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h1e == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_4(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h24 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_5(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h28 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_6(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h2e == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_7(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h32 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_8(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h38 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_9(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h3c == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_10(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h42 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_11(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h46 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_12(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h4c == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_13(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h50 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_14(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h56 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_15(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h5a == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_16(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h60 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_17(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h64 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_18(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h6a == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_19(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h6e == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_20(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h74 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_21(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h78 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_22(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h7e == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_23(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h82 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_24(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h88 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_25(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h8c == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_26(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h92 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_27(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h96 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_28(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'h9c == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_29(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'ha0 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_30(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'ha6 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_31(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'haa == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_32(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hb0 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_33(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hb4 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_34(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hba == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_35(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hbe == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_36(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hc4 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module LSU_37(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_read_addr,
  input         io_hostInterface_read_data_ready,
  output        io_hostInterface_read_data_valid,
  output [31:0] io_hostInterface_read_data_bits,
  input  [5:0]  io_hostInterface_write_addr,
  output        io_hostInterface_write_data_ready,
  input         io_hostInterface_write_data_valid,
  input  [31:0] io_hostInterface_write_data_bits,
  input         io_hostInterface_cycle,
  input         io_en,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  output [31:0] io_out_0
);
  wire  Muxn_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_io_out; // @[LSU.scala 61:34]
  wire  Muxn_1_io_config; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_0; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_in_1; // @[LSU.scala 61:34]
  wire [31:0] Muxn_1_io_out; // @[LSU.scala 61:34]
  wire  DelayPipe_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_io_out; // @[LSU.scala 62:42]
  wire  DelayPipe_1_clock; // @[LSU.scala 62:42]
  wire  DelayPipe_1_reset; // @[LSU.scala 62:42]
  wire  DelayPipe_1_io_en; // @[LSU.scala 62:42]
  wire [2:0] DelayPipe_1_io_config; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_in; // @[LSU.scala 62:42]
  wire [31:0] DelayPipe_1_io_out; // @[LSU.scala 62:42]
  wire  mem_clock; // @[LSU.scala 83:19]
  wire  mem_io_enable; // @[LSU.scala 83:19]
  wire  mem_io_write_enable; // @[LSU.scala 83:19]
  wire [5:0] mem_io_addr; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataIn; // @[LSU.scala 83:19]
  wire [31:0] mem_io_dataOut; // @[LSU.scala 83:19]
  wire  cfg_clock; // @[LSU.scala 134:19]
  wire  cfg_reset; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_en; // @[LSU.scala 134:19]
  wire  cfg_io_cfg_addr; // @[LSU.scala 134:19]
  wire [31:0] cfg_io_cfg_data; // @[LSU.scala 134:19]
  wire [40:0] cfg_io_out_0; // @[LSU.scala 134:19]
  wire [7:0] cfg_base_addr = 7'h0 * 7'h40; // @[LSU.scala 74:33]
  wire [6:0] _GEN_11 = {{6'd0}, io_hostInterface_cycle}; // @[LSU.scala 79:47]
  wire [7:0] host_base_addr = _GEN_11 * 7'h40; // @[LSU.scala 79:47]
  wire [31:0] Oprand_0 = DelayPipe_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_12 = {{2'd0}, io_hostInterface_read_addr}; // @[LSU.scala 104:72]
  wire [7:0] _T_3 = _GEN_12 + host_base_addr; // @[LSU.scala 104:72]
  wire [7:0] _GEN_13 = {{2'd0}, io_hostInterface_write_addr}; // @[LSU.scala 108:73]
  wire [7:0] _T_6 = _GEN_13 + host_base_addr; // @[LSU.scala 108:73]
  wire [31:0] opmode = {{31'd0}, cfg_io_out_0[40]}; // @[LSU.scala 56:20 LSU.scala 167:9]
  wire  _T_7 = opmode == 32'h0; // @[LSU.scala 110:17]
  wire  _T_8 = ~io_en; // @[LSU.scala 112:23]
  wire [7:0] _GEN_14 = {{2'd0}, Oprand_0[5:0]}; // @[LSU.scala 113:57]
  wire [7:0] _T_11 = _GEN_14 + cfg_base_addr; // @[LSU.scala 113:57]
  wire  _T_12 = opmode == 32'h1; // @[LSU.scala 114:23]
  wire [31:0] Oprand_1 = DelayPipe_1_io_out; // @[LSU.scala 55:20 LSU.scala 71:17]
  wire [7:0] _GEN_15 = {{2'd0}, Oprand_1[5:0]}; // @[LSU.scala 117:57]
  wire [7:0] _T_15 = _GEN_15 + cfg_base_addr; // @[LSU.scala 117:57]
  wire  _GEN_0 = _T_12 & io_en; // @[LSU.scala 114:32]
  wire [7:0] _GEN_1 = _T_12 ? _T_15 : 8'h0; // @[LSU.scala 114:32]
  wire  _GEN_2 = _T_7 ? io_en : _GEN_0; // @[LSU.scala 110:26]
  wire  _GEN_3 = _T_7 ? _T_8 : _GEN_0; // @[LSU.scala 110:26]
  wire [7:0] _GEN_4 = _T_7 ? _T_11 : _GEN_1; // @[LSU.scala 110:26]
  wire  _GEN_5 = io_hostInterface_write_data_valid | _GEN_2; // @[LSU.scala 105:49]
  wire  _GEN_6 = io_hostInterface_write_data_valid | _GEN_3; // @[LSU.scala 105:49]
  wire [7:0] _GEN_7 = io_hostInterface_write_data_valid ? _T_6 : _GEN_4; // @[LSU.scala 105:49]
  wire [7:0] _GEN_10 = io_hostInterface_read_data_ready ? _T_3 : _GEN_7; // @[LSU.scala 101:42]
  wire  _T_17 = 10'hc8 == io_cfg_addr[13:4]; // @[LSU.scala 135:48]
  wire [40:0] cfgOut = cfg_io_out_0; // @[LSU.scala 148:20 LSU.scala 149:10]
  Muxn Muxn ( // @[LSU.scala 61:34]
    .io_config(Muxn_io_config),
    .io_in_0(Muxn_io_in_0),
    .io_in_1(Muxn_io_in_1),
    .io_out(Muxn_io_out)
  );
  Muxn Muxn_1 ( // @[LSU.scala 61:34]
    .io_config(Muxn_1_io_config),
    .io_in_0(Muxn_1_io_in_0),
    .io_in_1(Muxn_1_io_in_1),
    .io_out(Muxn_1_io_out)
  );
  DelayPipe DelayPipe ( // @[LSU.scala 62:42]
    .clock(DelayPipe_clock),
    .reset(DelayPipe_reset),
    .io_en(DelayPipe_io_en),
    .io_config(DelayPipe_io_config),
    .io_in(DelayPipe_io_in),
    .io_out(DelayPipe_io_out)
  );
  DelayPipe DelayPipe_1 ( // @[LSU.scala 62:42]
    .clock(DelayPipe_1_clock),
    .reset(DelayPipe_1_reset),
    .io_en(DelayPipe_1_io_en),
    .io_config(DelayPipe_1_io_config),
    .io_in(DelayPipe_1_io_in),
    .io_out(DelayPipe_1_io_out)
  );
  single_port_ram mem ( // @[LSU.scala 83:19]
    .clock(mem_clock),
    .io_enable(mem_io_enable),
    .io_write_enable(mem_io_write_enable),
    .io_addr(mem_io_addr),
    .io_dataIn(mem_io_dataIn),
    .io_dataOut(mem_io_dataOut)
  );
  ConfigMem_143 cfg ( // @[LSU.scala 134:19]
    .clock(cfg_clock),
    .reset(cfg_reset),
    .io_cfg_en(cfg_io_cfg_en),
    .io_cfg_addr(cfg_io_cfg_addr),
    .io_cfg_data(cfg_io_cfg_data),
    .io_out_0(cfg_io_out_0)
  );
  assign io_hostInterface_read_data_valid = io_hostInterface_read_data_ready; // @[LSU.scala 93:36]
  assign io_hostInterface_read_data_bits = mem_io_dataOut; // @[LSU.scala 91:35]
  assign io_hostInterface_write_data_ready = io_hostInterface_write_data_valid; // @[LSU.scala 96:37]
  assign io_out_0 = mem_io_dataOut; // @[LSU.scala 87:13]
  assign Muxn_io_config = cfgOut[32]; // @[LSU.scala 154:20]
  assign Muxn_io_in_0 = io_in_0; // @[LSU.scala 66:23]
  assign Muxn_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign Muxn_1_io_config = cfgOut[33]; // @[LSU.scala 154:20]
  assign Muxn_1_io_in_0 = io_in_1; // @[LSU.scala 66:23]
  assign Muxn_1_io_in_1 = cfgOut[31:0]; // @[LSU.scala 68:29]
  assign DelayPipe_clock = clock;
  assign DelayPipe_reset = reset;
  assign DelayPipe_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_io_config = cfgOut[36:34]; // @[LSU.scala 160:29]
  assign DelayPipe_io_in = Muxn_io_out; // @[LSU.scala 70:25]
  assign DelayPipe_1_clock = clock;
  assign DelayPipe_1_reset = reset;
  assign DelayPipe_1_io_en = io_en; // @[LSU.scala 69:25]
  assign DelayPipe_1_io_config = cfgOut[39:37]; // @[LSU.scala 160:29]
  assign DelayPipe_1_io_in = Muxn_1_io_out; // @[LSU.scala 70:25]
  assign mem_clock = clock;
  assign mem_io_enable = io_hostInterface_read_data_ready | _GEN_5; // @[LSU.scala 84:17]
  assign mem_io_write_enable = io_hostInterface_read_data_ready ? 1'h0 : _GEN_6; // @[LSU.scala 85:23]
  assign mem_io_addr = _GEN_10[5:0]; // @[LSU.scala 86:15]
  assign mem_io_dataIn = io_hostInterface_write_data_valid ? io_hostInterface_write_data_bits : Oprand_0; // @[LSU.scala 88:17]
  assign cfg_clock = clock;
  assign cfg_reset = reset;
  assign cfg_io_cfg_en = io_cfg_en & _T_17; // @[LSU.scala 135:17]
  assign cfg_io_cfg_addr = io_cfg_addr[2]; // @[LSU.scala 136:19]
  assign cfg_io_cfg_data = io_cfg_data; // @[LSU.scala 140:19]
endmodule
module CGRA(
  input         clock,
  input         reset,
  input         io_cfg_en,
  input  [13:0] io_cfg_addr,
  input  [31:0] io_cfg_data,
  input  [5:0]  io_hostInterface_0_read_addr,
  input         io_hostInterface_0_read_data_ready,
  output        io_hostInterface_0_read_data_valid,
  output [31:0] io_hostInterface_0_read_data_bits,
  input  [5:0]  io_hostInterface_0_write_addr,
  output        io_hostInterface_0_write_data_ready,
  input         io_hostInterface_0_write_data_valid,
  input  [31:0] io_hostInterface_0_write_data_bits,
  input         io_hostInterface_0_cycle,
  input  [5:0]  io_hostInterface_1_read_addr,
  input         io_hostInterface_1_read_data_ready,
  output        io_hostInterface_1_read_data_valid,
  output [31:0] io_hostInterface_1_read_data_bits,
  input  [5:0]  io_hostInterface_1_write_addr,
  output        io_hostInterface_1_write_data_ready,
  input         io_hostInterface_1_write_data_valid,
  input  [31:0] io_hostInterface_1_write_data_bits,
  input         io_hostInterface_1_cycle,
  input  [5:0]  io_hostInterface_2_read_addr,
  input         io_hostInterface_2_read_data_ready,
  output        io_hostInterface_2_read_data_valid,
  output [31:0] io_hostInterface_2_read_data_bits,
  input  [5:0]  io_hostInterface_2_write_addr,
  output        io_hostInterface_2_write_data_ready,
  input         io_hostInterface_2_write_data_valid,
  input  [31:0] io_hostInterface_2_write_data_bits,
  input         io_hostInterface_2_cycle,
  input  [5:0]  io_hostInterface_3_read_addr,
  input         io_hostInterface_3_read_data_ready,
  output        io_hostInterface_3_read_data_valid,
  output [31:0] io_hostInterface_3_read_data_bits,
  input  [5:0]  io_hostInterface_3_write_addr,
  output        io_hostInterface_3_write_data_ready,
  input         io_hostInterface_3_write_data_valid,
  input  [31:0] io_hostInterface_3_write_data_bits,
  input         io_hostInterface_3_cycle,
  input  [5:0]  io_hostInterface_4_read_addr,
  input         io_hostInterface_4_read_data_ready,
  output        io_hostInterface_4_read_data_valid,
  output [31:0] io_hostInterface_4_read_data_bits,
  input  [5:0]  io_hostInterface_4_write_addr,
  output        io_hostInterface_4_write_data_ready,
  input         io_hostInterface_4_write_data_valid,
  input  [31:0] io_hostInterface_4_write_data_bits,
  input         io_hostInterface_4_cycle,
  input  [5:0]  io_hostInterface_5_read_addr,
  input         io_hostInterface_5_read_data_ready,
  output        io_hostInterface_5_read_data_valid,
  output [31:0] io_hostInterface_5_read_data_bits,
  input  [5:0]  io_hostInterface_5_write_addr,
  output        io_hostInterface_5_write_data_ready,
  input         io_hostInterface_5_write_data_valid,
  input  [31:0] io_hostInterface_5_write_data_bits,
  input         io_hostInterface_5_cycle,
  input  [5:0]  io_hostInterface_6_read_addr,
  input         io_hostInterface_6_read_data_ready,
  output        io_hostInterface_6_read_data_valid,
  output [31:0] io_hostInterface_6_read_data_bits,
  input  [5:0]  io_hostInterface_6_write_addr,
  output        io_hostInterface_6_write_data_ready,
  input         io_hostInterface_6_write_data_valid,
  input  [31:0] io_hostInterface_6_write_data_bits,
  input         io_hostInterface_6_cycle,
  input  [5:0]  io_hostInterface_7_read_addr,
  input         io_hostInterface_7_read_data_ready,
  output        io_hostInterface_7_read_data_valid,
  output [31:0] io_hostInterface_7_read_data_bits,
  input  [5:0]  io_hostInterface_7_write_addr,
  output        io_hostInterface_7_write_data_ready,
  input         io_hostInterface_7_write_data_valid,
  input  [31:0] io_hostInterface_7_write_data_bits,
  input         io_hostInterface_7_cycle,
  input  [5:0]  io_hostInterface_8_read_addr,
  input         io_hostInterface_8_read_data_ready,
  output        io_hostInterface_8_read_data_valid,
  output [31:0] io_hostInterface_8_read_data_bits,
  input  [5:0]  io_hostInterface_8_write_addr,
  output        io_hostInterface_8_write_data_ready,
  input         io_hostInterface_8_write_data_valid,
  input  [31:0] io_hostInterface_8_write_data_bits,
  input         io_hostInterface_8_cycle,
  input  [5:0]  io_hostInterface_9_read_addr,
  input         io_hostInterface_9_read_data_ready,
  output        io_hostInterface_9_read_data_valid,
  output [31:0] io_hostInterface_9_read_data_bits,
  input  [5:0]  io_hostInterface_9_write_addr,
  output        io_hostInterface_9_write_data_ready,
  input         io_hostInterface_9_write_data_valid,
  input  [31:0] io_hostInterface_9_write_data_bits,
  input         io_hostInterface_9_cycle,
  input  [5:0]  io_hostInterface_10_read_addr,
  input         io_hostInterface_10_read_data_ready,
  output        io_hostInterface_10_read_data_valid,
  output [31:0] io_hostInterface_10_read_data_bits,
  input  [5:0]  io_hostInterface_10_write_addr,
  output        io_hostInterface_10_write_data_ready,
  input         io_hostInterface_10_write_data_valid,
  input  [31:0] io_hostInterface_10_write_data_bits,
  input         io_hostInterface_10_cycle,
  input  [5:0]  io_hostInterface_11_read_addr,
  input         io_hostInterface_11_read_data_ready,
  output        io_hostInterface_11_read_data_valid,
  output [31:0] io_hostInterface_11_read_data_bits,
  input  [5:0]  io_hostInterface_11_write_addr,
  output        io_hostInterface_11_write_data_ready,
  input         io_hostInterface_11_write_data_valid,
  input  [31:0] io_hostInterface_11_write_data_bits,
  input         io_hostInterface_11_cycle,
  input  [5:0]  io_hostInterface_12_read_addr,
  input         io_hostInterface_12_read_data_ready,
  output        io_hostInterface_12_read_data_valid,
  output [31:0] io_hostInterface_12_read_data_bits,
  input  [5:0]  io_hostInterface_12_write_addr,
  output        io_hostInterface_12_write_data_ready,
  input         io_hostInterface_12_write_data_valid,
  input  [31:0] io_hostInterface_12_write_data_bits,
  input         io_hostInterface_12_cycle,
  input  [5:0]  io_hostInterface_13_read_addr,
  input         io_hostInterface_13_read_data_ready,
  output        io_hostInterface_13_read_data_valid,
  output [31:0] io_hostInterface_13_read_data_bits,
  input  [5:0]  io_hostInterface_13_write_addr,
  output        io_hostInterface_13_write_data_ready,
  input         io_hostInterface_13_write_data_valid,
  input  [31:0] io_hostInterface_13_write_data_bits,
  input         io_hostInterface_13_cycle,
  input  [5:0]  io_hostInterface_14_read_addr,
  input         io_hostInterface_14_read_data_ready,
  output        io_hostInterface_14_read_data_valid,
  output [31:0] io_hostInterface_14_read_data_bits,
  input  [5:0]  io_hostInterface_14_write_addr,
  output        io_hostInterface_14_write_data_ready,
  input         io_hostInterface_14_write_data_valid,
  input  [31:0] io_hostInterface_14_write_data_bits,
  input         io_hostInterface_14_cycle,
  input  [5:0]  io_hostInterface_15_read_addr,
  input         io_hostInterface_15_read_data_ready,
  output        io_hostInterface_15_read_data_valid,
  output [31:0] io_hostInterface_15_read_data_bits,
  input  [5:0]  io_hostInterface_15_write_addr,
  output        io_hostInterface_15_write_data_ready,
  input         io_hostInterface_15_write_data_valid,
  input  [31:0] io_hostInterface_15_write_data_bits,
  input         io_hostInterface_15_cycle,
  input  [5:0]  io_hostInterface_16_read_addr,
  input         io_hostInterface_16_read_data_ready,
  output        io_hostInterface_16_read_data_valid,
  output [31:0] io_hostInterface_16_read_data_bits,
  input  [5:0]  io_hostInterface_16_write_addr,
  output        io_hostInterface_16_write_data_ready,
  input         io_hostInterface_16_write_data_valid,
  input  [31:0] io_hostInterface_16_write_data_bits,
  input         io_hostInterface_16_cycle,
  input  [5:0]  io_hostInterface_17_read_addr,
  input         io_hostInterface_17_read_data_ready,
  output        io_hostInterface_17_read_data_valid,
  output [31:0] io_hostInterface_17_read_data_bits,
  input  [5:0]  io_hostInterface_17_write_addr,
  output        io_hostInterface_17_write_data_ready,
  input         io_hostInterface_17_write_data_valid,
  input  [31:0] io_hostInterface_17_write_data_bits,
  input         io_hostInterface_17_cycle,
  input  [5:0]  io_hostInterface_18_read_addr,
  input         io_hostInterface_18_read_data_ready,
  output        io_hostInterface_18_read_data_valid,
  output [31:0] io_hostInterface_18_read_data_bits,
  input  [5:0]  io_hostInterface_18_write_addr,
  output        io_hostInterface_18_write_data_ready,
  input         io_hostInterface_18_write_data_valid,
  input  [31:0] io_hostInterface_18_write_data_bits,
  input         io_hostInterface_18_cycle,
  input  [5:0]  io_hostInterface_19_read_addr,
  input         io_hostInterface_19_read_data_ready,
  output        io_hostInterface_19_read_data_valid,
  output [31:0] io_hostInterface_19_read_data_bits,
  input  [5:0]  io_hostInterface_19_write_addr,
  output        io_hostInterface_19_write_data_ready,
  input         io_hostInterface_19_write_data_valid,
  input  [31:0] io_hostInterface_19_write_data_bits,
  input         io_hostInterface_19_cycle,
  input  [5:0]  io_hostInterface_20_read_addr,
  input         io_hostInterface_20_read_data_ready,
  output        io_hostInterface_20_read_data_valid,
  output [31:0] io_hostInterface_20_read_data_bits,
  input  [5:0]  io_hostInterface_20_write_addr,
  output        io_hostInterface_20_write_data_ready,
  input         io_hostInterface_20_write_data_valid,
  input  [31:0] io_hostInterface_20_write_data_bits,
  input         io_hostInterface_20_cycle,
  input  [5:0]  io_hostInterface_21_read_addr,
  input         io_hostInterface_21_read_data_ready,
  output        io_hostInterface_21_read_data_valid,
  output [31:0] io_hostInterface_21_read_data_bits,
  input  [5:0]  io_hostInterface_21_write_addr,
  output        io_hostInterface_21_write_data_ready,
  input         io_hostInterface_21_write_data_valid,
  input  [31:0] io_hostInterface_21_write_data_bits,
  input         io_hostInterface_21_cycle,
  input  [5:0]  io_hostInterface_22_read_addr,
  input         io_hostInterface_22_read_data_ready,
  output        io_hostInterface_22_read_data_valid,
  output [31:0] io_hostInterface_22_read_data_bits,
  input  [5:0]  io_hostInterface_22_write_addr,
  output        io_hostInterface_22_write_data_ready,
  input         io_hostInterface_22_write_data_valid,
  input  [31:0] io_hostInterface_22_write_data_bits,
  input         io_hostInterface_22_cycle,
  input  [5:0]  io_hostInterface_23_read_addr,
  input         io_hostInterface_23_read_data_ready,
  output        io_hostInterface_23_read_data_valid,
  output [31:0] io_hostInterface_23_read_data_bits,
  input  [5:0]  io_hostInterface_23_write_addr,
  output        io_hostInterface_23_write_data_ready,
  input         io_hostInterface_23_write_data_valid,
  input  [31:0] io_hostInterface_23_write_data_bits,
  input         io_hostInterface_23_cycle,
  input  [5:0]  io_hostInterface_24_read_addr,
  input         io_hostInterface_24_read_data_ready,
  output        io_hostInterface_24_read_data_valid,
  output [31:0] io_hostInterface_24_read_data_bits,
  input  [5:0]  io_hostInterface_24_write_addr,
  output        io_hostInterface_24_write_data_ready,
  input         io_hostInterface_24_write_data_valid,
  input  [31:0] io_hostInterface_24_write_data_bits,
  input         io_hostInterface_24_cycle,
  input  [5:0]  io_hostInterface_25_read_addr,
  input         io_hostInterface_25_read_data_ready,
  output        io_hostInterface_25_read_data_valid,
  output [31:0] io_hostInterface_25_read_data_bits,
  input  [5:0]  io_hostInterface_25_write_addr,
  output        io_hostInterface_25_write_data_ready,
  input         io_hostInterface_25_write_data_valid,
  input  [31:0] io_hostInterface_25_write_data_bits,
  input         io_hostInterface_25_cycle,
  input  [5:0]  io_hostInterface_26_read_addr,
  input         io_hostInterface_26_read_data_ready,
  output        io_hostInterface_26_read_data_valid,
  output [31:0] io_hostInterface_26_read_data_bits,
  input  [5:0]  io_hostInterface_26_write_addr,
  output        io_hostInterface_26_write_data_ready,
  input         io_hostInterface_26_write_data_valid,
  input  [31:0] io_hostInterface_26_write_data_bits,
  input         io_hostInterface_26_cycle,
  input  [5:0]  io_hostInterface_27_read_addr,
  input         io_hostInterface_27_read_data_ready,
  output        io_hostInterface_27_read_data_valid,
  output [31:0] io_hostInterface_27_read_data_bits,
  input  [5:0]  io_hostInterface_27_write_addr,
  output        io_hostInterface_27_write_data_ready,
  input         io_hostInterface_27_write_data_valid,
  input  [31:0] io_hostInterface_27_write_data_bits,
  input         io_hostInterface_27_cycle,
  input  [5:0]  io_hostInterface_28_read_addr,
  input         io_hostInterface_28_read_data_ready,
  output        io_hostInterface_28_read_data_valid,
  output [31:0] io_hostInterface_28_read_data_bits,
  input  [5:0]  io_hostInterface_28_write_addr,
  output        io_hostInterface_28_write_data_ready,
  input         io_hostInterface_28_write_data_valid,
  input  [31:0] io_hostInterface_28_write_data_bits,
  input         io_hostInterface_28_cycle,
  input  [5:0]  io_hostInterface_29_read_addr,
  input         io_hostInterface_29_read_data_ready,
  output        io_hostInterface_29_read_data_valid,
  output [31:0] io_hostInterface_29_read_data_bits,
  input  [5:0]  io_hostInterface_29_write_addr,
  output        io_hostInterface_29_write_data_ready,
  input         io_hostInterface_29_write_data_valid,
  input  [31:0] io_hostInterface_29_write_data_bits,
  input         io_hostInterface_29_cycle,
  input  [5:0]  io_hostInterface_30_read_addr,
  input         io_hostInterface_30_read_data_ready,
  output        io_hostInterface_30_read_data_valid,
  output [31:0] io_hostInterface_30_read_data_bits,
  input  [5:0]  io_hostInterface_30_write_addr,
  output        io_hostInterface_30_write_data_ready,
  input         io_hostInterface_30_write_data_valid,
  input  [31:0] io_hostInterface_30_write_data_bits,
  input         io_hostInterface_30_cycle,
  input  [5:0]  io_hostInterface_31_read_addr,
  input         io_hostInterface_31_read_data_ready,
  output        io_hostInterface_31_read_data_valid,
  output [31:0] io_hostInterface_31_read_data_bits,
  input  [5:0]  io_hostInterface_31_write_addr,
  output        io_hostInterface_31_write_data_ready,
  input         io_hostInterface_31_write_data_valid,
  input  [31:0] io_hostInterface_31_write_data_bits,
  input         io_hostInterface_31_cycle,
  input  [5:0]  io_hostInterface_32_read_addr,
  input         io_hostInterface_32_read_data_ready,
  output        io_hostInterface_32_read_data_valid,
  output [31:0] io_hostInterface_32_read_data_bits,
  input  [5:0]  io_hostInterface_32_write_addr,
  output        io_hostInterface_32_write_data_ready,
  input         io_hostInterface_32_write_data_valid,
  input  [31:0] io_hostInterface_32_write_data_bits,
  input         io_hostInterface_32_cycle,
  input  [5:0]  io_hostInterface_33_read_addr,
  input         io_hostInterface_33_read_data_ready,
  output        io_hostInterface_33_read_data_valid,
  output [31:0] io_hostInterface_33_read_data_bits,
  input  [5:0]  io_hostInterface_33_write_addr,
  output        io_hostInterface_33_write_data_ready,
  input         io_hostInterface_33_write_data_valid,
  input  [31:0] io_hostInterface_33_write_data_bits,
  input         io_hostInterface_33_cycle,
  input  [5:0]  io_hostInterface_34_read_addr,
  input         io_hostInterface_34_read_data_ready,
  output        io_hostInterface_34_read_data_valid,
  output [31:0] io_hostInterface_34_read_data_bits,
  input  [5:0]  io_hostInterface_34_write_addr,
  output        io_hostInterface_34_write_data_ready,
  input         io_hostInterface_34_write_data_valid,
  input  [31:0] io_hostInterface_34_write_data_bits,
  input         io_hostInterface_34_cycle,
  input  [5:0]  io_hostInterface_35_read_addr,
  input         io_hostInterface_35_read_data_ready,
  output        io_hostInterface_35_read_data_valid,
  output [31:0] io_hostInterface_35_read_data_bits,
  input  [5:0]  io_hostInterface_35_write_addr,
  output        io_hostInterface_35_write_data_ready,
  input         io_hostInterface_35_write_data_valid,
  input  [31:0] io_hostInterface_35_write_data_bits,
  input         io_hostInterface_35_cycle,
  input  [5:0]  io_hostInterface_36_read_addr,
  input         io_hostInterface_36_read_data_ready,
  output        io_hostInterface_36_read_data_valid,
  output [31:0] io_hostInterface_36_read_data_bits,
  input  [5:0]  io_hostInterface_36_write_addr,
  output        io_hostInterface_36_write_data_ready,
  input         io_hostInterface_36_write_data_valid,
  input  [31:0] io_hostInterface_36_write_data_bits,
  input         io_hostInterface_36_cycle,
  input  [5:0]  io_hostInterface_37_read_addr,
  input         io_hostInterface_37_read_data_ready,
  output        io_hostInterface_37_read_data_valid,
  output [31:0] io_hostInterface_37_read_data_bits,
  input  [5:0]  io_hostInterface_37_write_addr,
  output        io_hostInterface_37_write_data_ready,
  input         io_hostInterface_37_write_data_valid,
  input  [31:0] io_hostInterface_37_write_data_bits,
  input         io_hostInterface_37_cycle,
  input         io_en_0,
  input         io_en_1,
  input         io_en_2,
  input         io_en_3,
  input         io_en_4,
  input  [31:0] io_in_0,
  input  [31:0] io_in_1,
  input  [31:0] io_in_2,
  input  [31:0] io_in_3,
  input  [31:0] io_in_4,
  input  [31:0] io_in_5,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3,
  output [31:0] io_out_4,
  output [31:0] io_out_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] ibs_0_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_0_io_out_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_1_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_1_io_out_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_2_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_2_io_out_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_3_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_3_io_out_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_4_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_4_io_out_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_5_io_in_0; // @[CGRA.scala 189:20]
  wire [31:0] ibs_5_io_out_0; // @[CGRA.scala 189:20]
  wire  obs_0_clock; // @[CGRA.scala 217:20]
  wire  obs_0_reset; // @[CGRA.scala 217:20]
  wire  obs_0_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_0_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_0_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_0_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_0_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_0_io_out_0; // @[CGRA.scala 217:20]
  wire  obs_1_clock; // @[CGRA.scala 217:20]
  wire  obs_1_reset; // @[CGRA.scala 217:20]
  wire  obs_1_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_1_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_1_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_1_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_1_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_1_io_out_0; // @[CGRA.scala 217:20]
  wire  obs_2_clock; // @[CGRA.scala 217:20]
  wire  obs_2_reset; // @[CGRA.scala 217:20]
  wire  obs_2_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_2_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_2_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_2_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_2_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_2_io_out_0; // @[CGRA.scala 217:20]
  wire  obs_3_clock; // @[CGRA.scala 217:20]
  wire  obs_3_reset; // @[CGRA.scala 217:20]
  wire  obs_3_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_3_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_3_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_3_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_3_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_3_io_out_0; // @[CGRA.scala 217:20]
  wire  obs_4_clock; // @[CGRA.scala 217:20]
  wire  obs_4_reset; // @[CGRA.scala 217:20]
  wire  obs_4_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_4_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_4_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_4_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_4_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_4_io_out_0; // @[CGRA.scala 217:20]
  wire  obs_5_clock; // @[CGRA.scala 217:20]
  wire  obs_5_reset; // @[CGRA.scala 217:20]
  wire  obs_5_io_cfg_en; // @[CGRA.scala 217:20]
  wire [13:0] obs_5_io_cfg_addr; // @[CGRA.scala 217:20]
  wire [31:0] obs_5_io_cfg_data; // @[CGRA.scala 217:20]
  wire [31:0] obs_5_io_in_0; // @[CGRA.scala 217:20]
  wire [31:0] obs_5_io_in_1; // @[CGRA.scala 217:20]
  wire [31:0] obs_5_io_out_0; // @[CGRA.scala 217:20]
  wire  pes_0_clock; // @[CGRA.scala 242:20]
  wire  pes_0_reset; // @[CGRA.scala 242:20]
  wire  pes_0_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_0_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_0_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_0_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_1_clock; // @[CGRA.scala 242:20]
  wire  pes_1_reset; // @[CGRA.scala 242:20]
  wire  pes_1_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_1_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_1_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_1_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_2_clock; // @[CGRA.scala 242:20]
  wire  pes_2_reset; // @[CGRA.scala 242:20]
  wire  pes_2_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_2_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_2_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_2_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_3_clock; // @[CGRA.scala 242:20]
  wire  pes_3_reset; // @[CGRA.scala 242:20]
  wire  pes_3_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_3_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_3_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_3_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_4_clock; // @[CGRA.scala 242:20]
  wire  pes_4_reset; // @[CGRA.scala 242:20]
  wire  pes_4_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_4_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_4_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_4_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_5_clock; // @[CGRA.scala 242:20]
  wire  pes_5_reset; // @[CGRA.scala 242:20]
  wire  pes_5_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_5_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_5_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_5_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_6_clock; // @[CGRA.scala 242:20]
  wire  pes_6_reset; // @[CGRA.scala 242:20]
  wire  pes_6_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_6_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_6_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_6_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_7_clock; // @[CGRA.scala 242:20]
  wire  pes_7_reset; // @[CGRA.scala 242:20]
  wire  pes_7_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_7_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_7_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_7_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_8_clock; // @[CGRA.scala 242:20]
  wire  pes_8_reset; // @[CGRA.scala 242:20]
  wire  pes_8_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_8_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_8_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_8_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_9_clock; // @[CGRA.scala 242:20]
  wire  pes_9_reset; // @[CGRA.scala 242:20]
  wire  pes_9_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_9_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_9_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_9_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_10_clock; // @[CGRA.scala 242:20]
  wire  pes_10_reset; // @[CGRA.scala 242:20]
  wire  pes_10_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_10_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_10_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_10_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_11_clock; // @[CGRA.scala 242:20]
  wire  pes_11_reset; // @[CGRA.scala 242:20]
  wire  pes_11_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_11_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_11_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_11_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_12_clock; // @[CGRA.scala 242:20]
  wire  pes_12_reset; // @[CGRA.scala 242:20]
  wire  pes_12_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_12_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_12_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_12_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_13_clock; // @[CGRA.scala 242:20]
  wire  pes_13_reset; // @[CGRA.scala 242:20]
  wire  pes_13_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_13_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_13_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_13_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_14_clock; // @[CGRA.scala 242:20]
  wire  pes_14_reset; // @[CGRA.scala 242:20]
  wire  pes_14_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_14_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_14_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_14_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_15_clock; // @[CGRA.scala 242:20]
  wire  pes_15_reset; // @[CGRA.scala 242:20]
  wire  pes_15_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_15_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_15_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_15_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_16_clock; // @[CGRA.scala 242:20]
  wire  pes_16_reset; // @[CGRA.scala 242:20]
  wire  pes_16_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_16_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_16_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_16_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_17_clock; // @[CGRA.scala 242:20]
  wire  pes_17_reset; // @[CGRA.scala 242:20]
  wire  pes_17_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_17_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_17_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_17_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_18_clock; // @[CGRA.scala 242:20]
  wire  pes_18_reset; // @[CGRA.scala 242:20]
  wire  pes_18_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_18_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_18_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_18_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_19_clock; // @[CGRA.scala 242:20]
  wire  pes_19_reset; // @[CGRA.scala 242:20]
  wire  pes_19_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_19_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_19_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_19_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_20_clock; // @[CGRA.scala 242:20]
  wire  pes_20_reset; // @[CGRA.scala 242:20]
  wire  pes_20_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_20_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_20_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_20_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_21_clock; // @[CGRA.scala 242:20]
  wire  pes_21_reset; // @[CGRA.scala 242:20]
  wire  pes_21_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_21_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_21_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_21_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_22_clock; // @[CGRA.scala 242:20]
  wire  pes_22_reset; // @[CGRA.scala 242:20]
  wire  pes_22_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_22_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_22_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_22_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_23_clock; // @[CGRA.scala 242:20]
  wire  pes_23_reset; // @[CGRA.scala 242:20]
  wire  pes_23_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_23_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_23_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_23_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_24_clock; // @[CGRA.scala 242:20]
  wire  pes_24_reset; // @[CGRA.scala 242:20]
  wire  pes_24_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_24_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_24_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_24_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_25_clock; // @[CGRA.scala 242:20]
  wire  pes_25_reset; // @[CGRA.scala 242:20]
  wire  pes_25_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_25_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_25_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_25_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_26_clock; // @[CGRA.scala 242:20]
  wire  pes_26_reset; // @[CGRA.scala 242:20]
  wire  pes_26_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_26_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_26_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_26_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_27_clock; // @[CGRA.scala 242:20]
  wire  pes_27_reset; // @[CGRA.scala 242:20]
  wire  pes_27_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_27_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_27_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_27_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_28_clock; // @[CGRA.scala 242:20]
  wire  pes_28_reset; // @[CGRA.scala 242:20]
  wire  pes_28_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_28_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_28_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_28_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_29_clock; // @[CGRA.scala 242:20]
  wire  pes_29_reset; // @[CGRA.scala 242:20]
  wire  pes_29_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_29_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_29_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_29_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_30_clock; // @[CGRA.scala 242:20]
  wire  pes_30_reset; // @[CGRA.scala 242:20]
  wire  pes_30_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_30_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_30_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_30_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_31_clock; // @[CGRA.scala 242:20]
  wire  pes_31_reset; // @[CGRA.scala 242:20]
  wire  pes_31_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_31_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_31_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_31_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_32_clock; // @[CGRA.scala 242:20]
  wire  pes_32_reset; // @[CGRA.scala 242:20]
  wire  pes_32_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_32_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_32_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_32_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_33_clock; // @[CGRA.scala 242:20]
  wire  pes_33_reset; // @[CGRA.scala 242:20]
  wire  pes_33_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_33_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_33_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_33_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_34_clock; // @[CGRA.scala 242:20]
  wire  pes_34_reset; // @[CGRA.scala 242:20]
  wire  pes_34_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_34_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_34_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_34_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_35_clock; // @[CGRA.scala 242:20]
  wire  pes_35_reset; // @[CGRA.scala 242:20]
  wire  pes_35_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_35_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_35_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_35_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_36_clock; // @[CGRA.scala 242:20]
  wire  pes_36_reset; // @[CGRA.scala 242:20]
  wire  pes_36_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_36_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_36_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_36_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_37_clock; // @[CGRA.scala 242:20]
  wire  pes_37_reset; // @[CGRA.scala 242:20]
  wire  pes_37_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_37_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_37_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_37_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_38_clock; // @[CGRA.scala 242:20]
  wire  pes_38_reset; // @[CGRA.scala 242:20]
  wire  pes_38_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_38_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_38_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_38_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_39_clock; // @[CGRA.scala 242:20]
  wire  pes_39_reset; // @[CGRA.scala 242:20]
  wire  pes_39_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_39_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_39_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_39_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_40_clock; // @[CGRA.scala 242:20]
  wire  pes_40_reset; // @[CGRA.scala 242:20]
  wire  pes_40_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_40_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_40_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_40_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_41_clock; // @[CGRA.scala 242:20]
  wire  pes_41_reset; // @[CGRA.scala 242:20]
  wire  pes_41_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_41_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_41_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_41_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_42_clock; // @[CGRA.scala 242:20]
  wire  pes_42_reset; // @[CGRA.scala 242:20]
  wire  pes_42_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_42_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_42_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_42_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_43_clock; // @[CGRA.scala 242:20]
  wire  pes_43_reset; // @[CGRA.scala 242:20]
  wire  pes_43_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_43_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_43_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_43_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_44_clock; // @[CGRA.scala 242:20]
  wire  pes_44_reset; // @[CGRA.scala 242:20]
  wire  pes_44_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_44_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_44_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_44_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_45_clock; // @[CGRA.scala 242:20]
  wire  pes_45_reset; // @[CGRA.scala 242:20]
  wire  pes_45_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_45_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_45_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_45_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_46_clock; // @[CGRA.scala 242:20]
  wire  pes_46_reset; // @[CGRA.scala 242:20]
  wire  pes_46_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_46_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_46_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_46_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_47_clock; // @[CGRA.scala 242:20]
  wire  pes_47_reset; // @[CGRA.scala 242:20]
  wire  pes_47_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_47_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_47_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_47_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_48_clock; // @[CGRA.scala 242:20]
  wire  pes_48_reset; // @[CGRA.scala 242:20]
  wire  pes_48_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_48_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_48_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_48_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_49_clock; // @[CGRA.scala 242:20]
  wire  pes_49_reset; // @[CGRA.scala 242:20]
  wire  pes_49_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_49_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_49_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_49_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_50_clock; // @[CGRA.scala 242:20]
  wire  pes_50_reset; // @[CGRA.scala 242:20]
  wire  pes_50_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_50_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_50_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_50_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_51_clock; // @[CGRA.scala 242:20]
  wire  pes_51_reset; // @[CGRA.scala 242:20]
  wire  pes_51_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_51_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_51_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_51_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_52_clock; // @[CGRA.scala 242:20]
  wire  pes_52_reset; // @[CGRA.scala 242:20]
  wire  pes_52_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_52_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_52_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_52_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_53_clock; // @[CGRA.scala 242:20]
  wire  pes_53_reset; // @[CGRA.scala 242:20]
  wire  pes_53_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_53_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_53_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_53_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_54_clock; // @[CGRA.scala 242:20]
  wire  pes_54_reset; // @[CGRA.scala 242:20]
  wire  pes_54_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_54_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_54_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_54_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_55_clock; // @[CGRA.scala 242:20]
  wire  pes_55_reset; // @[CGRA.scala 242:20]
  wire  pes_55_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_55_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_55_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_55_io_out_0; // @[CGRA.scala 242:20]
  wire  pes_56_clock; // @[CGRA.scala 242:20]
  wire  pes_56_reset; // @[CGRA.scala 242:20]
  wire  pes_56_io_cfg_en; // @[CGRA.scala 242:20]
  wire [13:0] pes_56_io_cfg_addr; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_cfg_data; // @[CGRA.scala 242:20]
  wire  pes_56_io_en; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_0; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_1; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_2; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_3; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_4; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_5; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_6; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_in_7; // @[CGRA.scala 242:20]
  wire [31:0] pes_56_io_out_0; // @[CGRA.scala 242:20]
  wire  gibs_0_clock; // @[CGRA.scala 333:21]
  wire  gibs_0_reset; // @[CGRA.scala 333:21]
  wire  gibs_0_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_0_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_0_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_1_clock; // @[CGRA.scala 333:21]
  wire  gibs_1_reset; // @[CGRA.scala 333:21]
  wire  gibs_1_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_1_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_1_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_2_clock; // @[CGRA.scala 333:21]
  wire  gibs_2_reset; // @[CGRA.scala 333:21]
  wire  gibs_2_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_2_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_2_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_3_clock; // @[CGRA.scala 333:21]
  wire  gibs_3_reset; // @[CGRA.scala 333:21]
  wire  gibs_3_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_3_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_3_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_4_clock; // @[CGRA.scala 333:21]
  wire  gibs_4_reset; // @[CGRA.scala 333:21]
  wire  gibs_4_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_4_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_4_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_5_clock; // @[CGRA.scala 333:21]
  wire  gibs_5_reset; // @[CGRA.scala 333:21]
  wire  gibs_5_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_5_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_5_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_6_clock; // @[CGRA.scala 333:21]
  wire  gibs_6_reset; // @[CGRA.scala 333:21]
  wire  gibs_6_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_6_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_6_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_7_clock; // @[CGRA.scala 333:21]
  wire  gibs_7_reset; // @[CGRA.scala 333:21]
  wire  gibs_7_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_7_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_7_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_8_clock; // @[CGRA.scala 333:21]
  wire  gibs_8_reset; // @[CGRA.scala 333:21]
  wire  gibs_8_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_8_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_8_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_9_clock; // @[CGRA.scala 333:21]
  wire  gibs_9_reset; // @[CGRA.scala 333:21]
  wire  gibs_9_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_9_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_9_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_10_clock; // @[CGRA.scala 333:21]
  wire  gibs_10_reset; // @[CGRA.scala 333:21]
  wire  gibs_10_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_10_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_10_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_11_clock; // @[CGRA.scala 333:21]
  wire  gibs_11_reset; // @[CGRA.scala 333:21]
  wire  gibs_11_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_11_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_11_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_12_clock; // @[CGRA.scala 333:21]
  wire  gibs_12_reset; // @[CGRA.scala 333:21]
  wire  gibs_12_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_12_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_12_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_13_clock; // @[CGRA.scala 333:21]
  wire  gibs_13_reset; // @[CGRA.scala 333:21]
  wire  gibs_13_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_13_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_13_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_14_clock; // @[CGRA.scala 333:21]
  wire  gibs_14_reset; // @[CGRA.scala 333:21]
  wire  gibs_14_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_14_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_14_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_15_clock; // @[CGRA.scala 333:21]
  wire  gibs_15_reset; // @[CGRA.scala 333:21]
  wire  gibs_15_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_15_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_15_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_16_clock; // @[CGRA.scala 333:21]
  wire  gibs_16_reset; // @[CGRA.scala 333:21]
  wire  gibs_16_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_16_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_16_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_17_clock; // @[CGRA.scala 333:21]
  wire  gibs_17_reset; // @[CGRA.scala 333:21]
  wire  gibs_17_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_17_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_17_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_18_clock; // @[CGRA.scala 333:21]
  wire  gibs_18_reset; // @[CGRA.scala 333:21]
  wire  gibs_18_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_18_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_18_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_19_clock; // @[CGRA.scala 333:21]
  wire  gibs_19_reset; // @[CGRA.scala 333:21]
  wire  gibs_19_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_19_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_19_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_20_clock; // @[CGRA.scala 333:21]
  wire  gibs_20_reset; // @[CGRA.scala 333:21]
  wire  gibs_20_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_20_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_20_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_21_clock; // @[CGRA.scala 333:21]
  wire  gibs_21_reset; // @[CGRA.scala 333:21]
  wire  gibs_21_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_21_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_21_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_22_clock; // @[CGRA.scala 333:21]
  wire  gibs_22_reset; // @[CGRA.scala 333:21]
  wire  gibs_22_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_22_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_22_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_23_clock; // @[CGRA.scala 333:21]
  wire  gibs_23_reset; // @[CGRA.scala 333:21]
  wire  gibs_23_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_23_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_23_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_24_clock; // @[CGRA.scala 333:21]
  wire  gibs_24_reset; // @[CGRA.scala 333:21]
  wire  gibs_24_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_24_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_24_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_25_clock; // @[CGRA.scala 333:21]
  wire  gibs_25_reset; // @[CGRA.scala 333:21]
  wire  gibs_25_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_25_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_25_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_26_clock; // @[CGRA.scala 333:21]
  wire  gibs_26_reset; // @[CGRA.scala 333:21]
  wire  gibs_26_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_26_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_26_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_27_clock; // @[CGRA.scala 333:21]
  wire  gibs_27_reset; // @[CGRA.scala 333:21]
  wire  gibs_27_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_27_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_27_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_28_clock; // @[CGRA.scala 333:21]
  wire  gibs_28_reset; // @[CGRA.scala 333:21]
  wire  gibs_28_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_28_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_28_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_29_clock; // @[CGRA.scala 333:21]
  wire  gibs_29_reset; // @[CGRA.scala 333:21]
  wire  gibs_29_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_29_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_29_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_30_clock; // @[CGRA.scala 333:21]
  wire  gibs_30_reset; // @[CGRA.scala 333:21]
  wire  gibs_30_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_30_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_30_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_31_clock; // @[CGRA.scala 333:21]
  wire  gibs_31_reset; // @[CGRA.scala 333:21]
  wire  gibs_31_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_31_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_31_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_32_clock; // @[CGRA.scala 333:21]
  wire  gibs_32_reset; // @[CGRA.scala 333:21]
  wire  gibs_32_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_32_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_32_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_33_clock; // @[CGRA.scala 333:21]
  wire  gibs_33_reset; // @[CGRA.scala 333:21]
  wire  gibs_33_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_33_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_33_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_34_clock; // @[CGRA.scala 333:21]
  wire  gibs_34_reset; // @[CGRA.scala 333:21]
  wire  gibs_34_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_34_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_34_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_35_clock; // @[CGRA.scala 333:21]
  wire  gibs_35_reset; // @[CGRA.scala 333:21]
  wire  gibs_35_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_35_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_35_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_36_clock; // @[CGRA.scala 333:21]
  wire  gibs_36_reset; // @[CGRA.scala 333:21]
  wire  gibs_36_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_36_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_36_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_37_clock; // @[CGRA.scala 333:21]
  wire  gibs_37_reset; // @[CGRA.scala 333:21]
  wire  gibs_37_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_37_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_37_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_38_clock; // @[CGRA.scala 333:21]
  wire  gibs_38_reset; // @[CGRA.scala 333:21]
  wire  gibs_38_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_38_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_38_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_39_clock; // @[CGRA.scala 333:21]
  wire  gibs_39_reset; // @[CGRA.scala 333:21]
  wire  gibs_39_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_39_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_39_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_40_clock; // @[CGRA.scala 333:21]
  wire  gibs_40_reset; // @[CGRA.scala 333:21]
  wire  gibs_40_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_40_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_40_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_41_clock; // @[CGRA.scala 333:21]
  wire  gibs_41_reset; // @[CGRA.scala 333:21]
  wire  gibs_41_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_41_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_41_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_42_clock; // @[CGRA.scala 333:21]
  wire  gibs_42_reset; // @[CGRA.scala 333:21]
  wire  gibs_42_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_42_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_42_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_43_clock; // @[CGRA.scala 333:21]
  wire  gibs_43_reset; // @[CGRA.scala 333:21]
  wire  gibs_43_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_43_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_43_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_44_clock; // @[CGRA.scala 333:21]
  wire  gibs_44_reset; // @[CGRA.scala 333:21]
  wire  gibs_44_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_44_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_44_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_45_clock; // @[CGRA.scala 333:21]
  wire  gibs_45_reset; // @[CGRA.scala 333:21]
  wire  gibs_45_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_45_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_45_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_46_clock; // @[CGRA.scala 333:21]
  wire  gibs_46_reset; // @[CGRA.scala 333:21]
  wire  gibs_46_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_46_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_46_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_47_clock; // @[CGRA.scala 333:21]
  wire  gibs_47_reset; // @[CGRA.scala 333:21]
  wire  gibs_47_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_47_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_47_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_48_clock; // @[CGRA.scala 333:21]
  wire  gibs_48_reset; // @[CGRA.scala 333:21]
  wire  gibs_48_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_48_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_48_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_49_clock; // @[CGRA.scala 333:21]
  wire  gibs_49_reset; // @[CGRA.scala 333:21]
  wire  gibs_49_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_49_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_49_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_50_clock; // @[CGRA.scala 333:21]
  wire  gibs_50_reset; // @[CGRA.scala 333:21]
  wire  gibs_50_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_50_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_50_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_51_clock; // @[CGRA.scala 333:21]
  wire  gibs_51_reset; // @[CGRA.scala 333:21]
  wire  gibs_51_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_51_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_51_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_52_clock; // @[CGRA.scala 333:21]
  wire  gibs_52_reset; // @[CGRA.scala 333:21]
  wire  gibs_52_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_52_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_52_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_53_clock; // @[CGRA.scala 333:21]
  wire  gibs_53_reset; // @[CGRA.scala 333:21]
  wire  gibs_53_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_53_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_53_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_54_clock; // @[CGRA.scala 333:21]
  wire  gibs_54_reset; // @[CGRA.scala 333:21]
  wire  gibs_54_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_54_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_54_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_55_clock; // @[CGRA.scala 333:21]
  wire  gibs_55_reset; // @[CGRA.scala 333:21]
  wire  gibs_55_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_55_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_55_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_56_clock; // @[CGRA.scala 333:21]
  wire  gibs_56_reset; // @[CGRA.scala 333:21]
  wire  gibs_56_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_56_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_56_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_57_clock; // @[CGRA.scala 333:21]
  wire  gibs_57_reset; // @[CGRA.scala 333:21]
  wire  gibs_57_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_57_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_57_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_58_clock; // @[CGRA.scala 333:21]
  wire  gibs_58_reset; // @[CGRA.scala 333:21]
  wire  gibs_58_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_58_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_58_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_59_clock; // @[CGRA.scala 333:21]
  wire  gibs_59_reset; // @[CGRA.scala 333:21]
  wire  gibs_59_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_59_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_59_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_60_clock; // @[CGRA.scala 333:21]
  wire  gibs_60_reset; // @[CGRA.scala 333:21]
  wire  gibs_60_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_60_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_60_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_61_clock; // @[CGRA.scala 333:21]
  wire  gibs_61_reset; // @[CGRA.scala 333:21]
  wire  gibs_61_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_61_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_61_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_62_clock; // @[CGRA.scala 333:21]
  wire  gibs_62_reset; // @[CGRA.scala 333:21]
  wire  gibs_62_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_62_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_62_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_63_clock; // @[CGRA.scala 333:21]
  wire  gibs_63_reset; // @[CGRA.scala 333:21]
  wire  gibs_63_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_63_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_63_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_64_clock; // @[CGRA.scala 333:21]
  wire  gibs_64_reset; // @[CGRA.scala 333:21]
  wire  gibs_64_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_64_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_64_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_65_clock; // @[CGRA.scala 333:21]
  wire  gibs_65_reset; // @[CGRA.scala 333:21]
  wire  gibs_65_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_65_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_65_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_66_clock; // @[CGRA.scala 333:21]
  wire  gibs_66_reset; // @[CGRA.scala 333:21]
  wire  gibs_66_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_66_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_66_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_67_clock; // @[CGRA.scala 333:21]
  wire  gibs_67_reset; // @[CGRA.scala 333:21]
  wire  gibs_67_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_67_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_67_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_68_clock; // @[CGRA.scala 333:21]
  wire  gibs_68_reset; // @[CGRA.scala 333:21]
  wire  gibs_68_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_68_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_68_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_69_clock; // @[CGRA.scala 333:21]
  wire  gibs_69_reset; // @[CGRA.scala 333:21]
  wire  gibs_69_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_69_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_69_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_70_clock; // @[CGRA.scala 333:21]
  wire  gibs_70_reset; // @[CGRA.scala 333:21]
  wire  gibs_70_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_70_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_70_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_71_clock; // @[CGRA.scala 333:21]
  wire  gibs_71_reset; // @[CGRA.scala 333:21]
  wire  gibs_71_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_71_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_71_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_72_clock; // @[CGRA.scala 333:21]
  wire  gibs_72_reset; // @[CGRA.scala 333:21]
  wire  gibs_72_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_72_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_72_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_73_clock; // @[CGRA.scala 333:21]
  wire  gibs_73_reset; // @[CGRA.scala 333:21]
  wire  gibs_73_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_73_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_73_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_74_clock; // @[CGRA.scala 333:21]
  wire  gibs_74_reset; // @[CGRA.scala 333:21]
  wire  gibs_74_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_74_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinSE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_otrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_74_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_75_clock; // @[CGRA.scala 333:21]
  wire  gibs_75_reset; // @[CGRA.scala 333:21]
  wire  gibs_75_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_75_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_ipinSW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_itrackS_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_75_io_otrackS_0; // @[CGRA.scala 333:21]
  wire  gibs_76_clock; // @[CGRA.scala 333:21]
  wire  gibs_76_reset; // @[CGRA.scala 333:21]
  wire  gibs_76_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_76_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_76_io_otrackE_0; // @[CGRA.scala 333:21]
  wire  gibs_77_clock; // @[CGRA.scala 333:21]
  wire  gibs_77_reset; // @[CGRA.scala 333:21]
  wire  gibs_77_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_77_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_77_io_otrackE_0; // @[CGRA.scala 333:21]
  wire  gibs_78_clock; // @[CGRA.scala 333:21]
  wire  gibs_78_reset; // @[CGRA.scala 333:21]
  wire  gibs_78_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_78_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinNE_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_opinSE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_otrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_itrackE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_78_io_otrackE_0; // @[CGRA.scala 333:21]
  wire  gibs_79_clock; // @[CGRA.scala 333:21]
  wire  gibs_79_reset; // @[CGRA.scala 333:21]
  wire  gibs_79_io_cfg_en; // @[CGRA.scala 333:21]
  wire [13:0] gibs_79_io_cfg_addr; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_cfg_data; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_ipinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_ipinNW_1; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_opinNW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_ipinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_opinNE_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_ipinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_opinSW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_itrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_otrackW_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_itrackN_0; // @[CGRA.scala 333:21]
  wire [31:0] gibs_79_io_otrackN_0; // @[CGRA.scala 333:21]
  wire  lsus_0_clock; // @[CGRA.scala 364:21]
  wire  lsus_0_reset; // @[CGRA.scala 364:21]
  wire  lsus_0_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_0_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_0_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_0_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_0_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_0_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_0_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_0_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_0_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_0_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_0_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_1_clock; // @[CGRA.scala 364:21]
  wire  lsus_1_reset; // @[CGRA.scala 364:21]
  wire  lsus_1_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_1_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_1_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_1_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_1_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_1_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_1_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_1_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_1_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_1_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_1_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_2_clock; // @[CGRA.scala 364:21]
  wire  lsus_2_reset; // @[CGRA.scala 364:21]
  wire  lsus_2_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_2_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_2_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_2_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_2_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_2_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_2_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_2_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_2_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_2_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_2_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_3_clock; // @[CGRA.scala 364:21]
  wire  lsus_3_reset; // @[CGRA.scala 364:21]
  wire  lsus_3_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_3_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_3_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_3_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_3_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_3_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_3_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_3_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_3_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_3_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_3_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_4_clock; // @[CGRA.scala 364:21]
  wire  lsus_4_reset; // @[CGRA.scala 364:21]
  wire  lsus_4_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_4_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_4_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_4_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_4_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_4_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_4_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_4_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_4_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_4_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_4_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_5_clock; // @[CGRA.scala 364:21]
  wire  lsus_5_reset; // @[CGRA.scala 364:21]
  wire  lsus_5_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_5_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_5_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_5_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_5_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_5_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_5_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_5_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_5_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_5_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_5_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_6_clock; // @[CGRA.scala 364:21]
  wire  lsus_6_reset; // @[CGRA.scala 364:21]
  wire  lsus_6_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_6_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_6_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_6_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_6_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_6_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_6_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_6_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_6_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_6_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_6_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_7_clock; // @[CGRA.scala 364:21]
  wire  lsus_7_reset; // @[CGRA.scala 364:21]
  wire  lsus_7_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_7_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_7_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_7_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_7_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_7_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_7_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_7_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_7_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_7_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_7_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_8_clock; // @[CGRA.scala 364:21]
  wire  lsus_8_reset; // @[CGRA.scala 364:21]
  wire  lsus_8_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_8_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_8_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_8_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_8_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_8_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_8_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_8_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_8_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_8_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_8_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_9_clock; // @[CGRA.scala 364:21]
  wire  lsus_9_reset; // @[CGRA.scala 364:21]
  wire  lsus_9_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_9_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_9_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_9_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_9_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_9_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_9_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_9_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_9_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_9_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_9_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_10_clock; // @[CGRA.scala 364:21]
  wire  lsus_10_reset; // @[CGRA.scala 364:21]
  wire  lsus_10_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_10_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_10_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_10_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_10_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_10_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_10_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_10_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_10_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_10_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_10_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_11_clock; // @[CGRA.scala 364:21]
  wire  lsus_11_reset; // @[CGRA.scala 364:21]
  wire  lsus_11_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_11_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_11_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_11_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_11_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_11_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_11_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_11_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_11_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_11_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_11_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_12_clock; // @[CGRA.scala 364:21]
  wire  lsus_12_reset; // @[CGRA.scala 364:21]
  wire  lsus_12_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_12_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_12_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_12_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_12_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_12_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_12_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_12_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_12_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_12_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_12_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_13_clock; // @[CGRA.scala 364:21]
  wire  lsus_13_reset; // @[CGRA.scala 364:21]
  wire  lsus_13_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_13_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_13_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_13_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_13_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_13_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_13_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_13_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_13_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_13_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_13_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_14_clock; // @[CGRA.scala 364:21]
  wire  lsus_14_reset; // @[CGRA.scala 364:21]
  wire  lsus_14_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_14_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_14_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_14_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_14_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_14_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_14_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_14_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_14_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_14_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_14_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_15_clock; // @[CGRA.scala 364:21]
  wire  lsus_15_reset; // @[CGRA.scala 364:21]
  wire  lsus_15_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_15_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_15_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_15_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_15_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_15_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_15_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_15_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_15_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_15_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_15_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_16_clock; // @[CGRA.scala 364:21]
  wire  lsus_16_reset; // @[CGRA.scala 364:21]
  wire  lsus_16_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_16_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_16_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_16_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_16_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_16_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_16_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_16_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_16_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_16_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_16_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_17_clock; // @[CGRA.scala 364:21]
  wire  lsus_17_reset; // @[CGRA.scala 364:21]
  wire  lsus_17_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_17_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_17_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_17_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_17_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_17_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_17_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_17_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_17_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_17_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_17_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_18_clock; // @[CGRA.scala 364:21]
  wire  lsus_18_reset; // @[CGRA.scala 364:21]
  wire  lsus_18_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_18_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_18_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_18_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_18_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_18_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_18_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_18_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_18_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_18_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_18_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_19_clock; // @[CGRA.scala 364:21]
  wire  lsus_19_reset; // @[CGRA.scala 364:21]
  wire  lsus_19_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_19_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_19_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_19_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_19_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_19_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_19_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_19_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_19_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_19_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_19_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_20_clock; // @[CGRA.scala 364:21]
  wire  lsus_20_reset; // @[CGRA.scala 364:21]
  wire  lsus_20_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_20_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_20_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_20_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_20_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_20_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_20_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_20_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_20_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_20_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_20_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_21_clock; // @[CGRA.scala 364:21]
  wire  lsus_21_reset; // @[CGRA.scala 364:21]
  wire  lsus_21_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_21_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_21_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_21_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_21_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_21_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_21_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_21_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_21_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_21_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_21_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_22_clock; // @[CGRA.scala 364:21]
  wire  lsus_22_reset; // @[CGRA.scala 364:21]
  wire  lsus_22_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_22_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_22_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_22_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_22_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_22_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_22_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_22_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_22_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_22_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_22_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_23_clock; // @[CGRA.scala 364:21]
  wire  lsus_23_reset; // @[CGRA.scala 364:21]
  wire  lsus_23_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_23_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_23_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_23_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_23_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_23_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_23_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_23_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_23_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_23_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_23_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_24_clock; // @[CGRA.scala 364:21]
  wire  lsus_24_reset; // @[CGRA.scala 364:21]
  wire  lsus_24_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_24_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_24_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_24_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_24_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_24_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_24_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_24_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_24_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_24_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_24_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_25_clock; // @[CGRA.scala 364:21]
  wire  lsus_25_reset; // @[CGRA.scala 364:21]
  wire  lsus_25_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_25_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_25_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_25_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_25_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_25_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_25_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_25_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_25_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_25_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_25_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_26_clock; // @[CGRA.scala 364:21]
  wire  lsus_26_reset; // @[CGRA.scala 364:21]
  wire  lsus_26_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_26_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_26_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_26_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_26_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_26_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_26_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_26_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_26_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_26_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_26_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_27_clock; // @[CGRA.scala 364:21]
  wire  lsus_27_reset; // @[CGRA.scala 364:21]
  wire  lsus_27_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_27_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_27_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_27_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_27_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_27_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_27_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_27_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_27_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_27_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_27_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_28_clock; // @[CGRA.scala 364:21]
  wire  lsus_28_reset; // @[CGRA.scala 364:21]
  wire  lsus_28_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_28_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_28_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_28_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_28_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_28_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_28_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_28_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_28_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_28_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_28_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_29_clock; // @[CGRA.scala 364:21]
  wire  lsus_29_reset; // @[CGRA.scala 364:21]
  wire  lsus_29_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_29_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_29_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_29_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_29_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_29_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_29_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_29_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_29_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_29_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_29_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_30_clock; // @[CGRA.scala 364:21]
  wire  lsus_30_reset; // @[CGRA.scala 364:21]
  wire  lsus_30_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_30_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_30_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_30_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_30_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_30_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_30_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_30_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_30_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_30_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_30_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_31_clock; // @[CGRA.scala 364:21]
  wire  lsus_31_reset; // @[CGRA.scala 364:21]
  wire  lsus_31_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_31_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_31_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_31_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_31_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_31_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_31_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_31_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_31_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_31_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_31_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_32_clock; // @[CGRA.scala 364:21]
  wire  lsus_32_reset; // @[CGRA.scala 364:21]
  wire  lsus_32_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_32_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_32_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_32_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_32_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_32_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_32_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_32_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_32_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_32_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_32_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_33_clock; // @[CGRA.scala 364:21]
  wire  lsus_33_reset; // @[CGRA.scala 364:21]
  wire  lsus_33_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_33_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_33_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_33_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_33_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_33_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_33_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_33_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_33_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_33_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_33_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_34_clock; // @[CGRA.scala 364:21]
  wire  lsus_34_reset; // @[CGRA.scala 364:21]
  wire  lsus_34_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_34_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_34_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_34_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_34_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_34_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_34_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_34_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_34_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_34_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_34_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_35_clock; // @[CGRA.scala 364:21]
  wire  lsus_35_reset; // @[CGRA.scala 364:21]
  wire  lsus_35_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_35_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_35_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_35_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_35_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_35_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_35_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_35_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_35_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_35_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_35_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_36_clock; // @[CGRA.scala 364:21]
  wire  lsus_36_reset; // @[CGRA.scala 364:21]
  wire  lsus_36_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_36_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_36_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_36_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_36_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_36_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_36_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_36_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_36_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_36_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_36_io_out_0; // @[CGRA.scala 364:21]
  wire  lsus_37_clock; // @[CGRA.scala 364:21]
  wire  lsus_37_reset; // @[CGRA.scala 364:21]
  wire  lsus_37_io_cfg_en; // @[CGRA.scala 364:21]
  wire [13:0] lsus_37_io_cfg_addr; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_cfg_data; // @[CGRA.scala 364:21]
  wire [5:0] lsus_37_io_hostInterface_read_addr; // @[CGRA.scala 364:21]
  wire  lsus_37_io_hostInterface_read_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_37_io_hostInterface_read_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_hostInterface_read_data_bits; // @[CGRA.scala 364:21]
  wire [5:0] lsus_37_io_hostInterface_write_addr; // @[CGRA.scala 364:21]
  wire  lsus_37_io_hostInterface_write_data_ready; // @[CGRA.scala 364:21]
  wire  lsus_37_io_hostInterface_write_data_valid; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_hostInterface_write_data_bits; // @[CGRA.scala 364:21]
  wire  lsus_37_io_hostInterface_cycle; // @[CGRA.scala 364:21]
  wire  lsus_37_io_en; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_in_0; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_in_1; // @[CGRA.scala 364:21]
  wire [31:0] lsus_37_io_out_0; // @[CGRA.scala 364:21]
  reg [46:0] cfgRegs_0; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_1; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_2; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_3; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_4; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_5; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_6; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_7; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_8; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_9; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_10; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_11; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_12; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_13; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_14; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_15; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_16; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_17; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_18; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_19; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_20; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_21; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_22; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_23; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_24; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_25; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_26; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_27; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_28; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_29; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_30; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_31; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_32; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_33; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_34; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_35; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_36; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_37; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_38; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_39; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_40; // @[CGRA.scala 645:24]
  reg [46:0] cfgRegs_41; // @[CGRA.scala 645:24]
  wire [46:0] _T_2 = {io_cfg_en,io_cfg_addr,io_cfg_data}; // @[Cat.scala 29:58]
  IOB ibs_0 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_0_io_in_0),
    .io_out_0(ibs_0_io_out_0)
  );
  IOB ibs_1 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_1_io_in_0),
    .io_out_0(ibs_1_io_out_0)
  );
  IOB ibs_2 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_2_io_in_0),
    .io_out_0(ibs_2_io_out_0)
  );
  IOB ibs_3 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_3_io_in_0),
    .io_out_0(ibs_3_io_out_0)
  );
  IOB ibs_4 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_4_io_in_0),
    .io_out_0(ibs_4_io_out_0)
  );
  IOB ibs_5 ( // @[CGRA.scala 189:20]
    .io_in_0(ibs_5_io_in_0),
    .io_out_0(ibs_5_io_out_0)
  );
  IOB_6 obs_0 ( // @[CGRA.scala 217:20]
    .clock(obs_0_clock),
    .reset(obs_0_reset),
    .io_cfg_en(obs_0_io_cfg_en),
    .io_cfg_addr(obs_0_io_cfg_addr),
    .io_cfg_data(obs_0_io_cfg_data),
    .io_in_0(obs_0_io_in_0),
    .io_in_1(obs_0_io_in_1),
    .io_out_0(obs_0_io_out_0)
  );
  IOB_7 obs_1 ( // @[CGRA.scala 217:20]
    .clock(obs_1_clock),
    .reset(obs_1_reset),
    .io_cfg_en(obs_1_io_cfg_en),
    .io_cfg_addr(obs_1_io_cfg_addr),
    .io_cfg_data(obs_1_io_cfg_data),
    .io_in_0(obs_1_io_in_0),
    .io_in_1(obs_1_io_in_1),
    .io_out_0(obs_1_io_out_0)
  );
  IOB_8 obs_2 ( // @[CGRA.scala 217:20]
    .clock(obs_2_clock),
    .reset(obs_2_reset),
    .io_cfg_en(obs_2_io_cfg_en),
    .io_cfg_addr(obs_2_io_cfg_addr),
    .io_cfg_data(obs_2_io_cfg_data),
    .io_in_0(obs_2_io_in_0),
    .io_in_1(obs_2_io_in_1),
    .io_out_0(obs_2_io_out_0)
  );
  IOB_9 obs_3 ( // @[CGRA.scala 217:20]
    .clock(obs_3_clock),
    .reset(obs_3_reset),
    .io_cfg_en(obs_3_io_cfg_en),
    .io_cfg_addr(obs_3_io_cfg_addr),
    .io_cfg_data(obs_3_io_cfg_data),
    .io_in_0(obs_3_io_in_0),
    .io_in_1(obs_3_io_in_1),
    .io_out_0(obs_3_io_out_0)
  );
  IOB_10 obs_4 ( // @[CGRA.scala 217:20]
    .clock(obs_4_clock),
    .reset(obs_4_reset),
    .io_cfg_en(obs_4_io_cfg_en),
    .io_cfg_addr(obs_4_io_cfg_addr),
    .io_cfg_data(obs_4_io_cfg_data),
    .io_in_0(obs_4_io_in_0),
    .io_in_1(obs_4_io_in_1),
    .io_out_0(obs_4_io_out_0)
  );
  IOB_11 obs_5 ( // @[CGRA.scala 217:20]
    .clock(obs_5_clock),
    .reset(obs_5_reset),
    .io_cfg_en(obs_5_io_cfg_en),
    .io_cfg_addr(obs_5_io_cfg_addr),
    .io_cfg_data(obs_5_io_cfg_data),
    .io_in_0(obs_5_io_in_0),
    .io_in_1(obs_5_io_in_1),
    .io_out_0(obs_5_io_out_0)
  );
  GPE pes_0 ( // @[CGRA.scala 242:20]
    .clock(pes_0_clock),
    .reset(pes_0_reset),
    .io_cfg_en(pes_0_io_cfg_en),
    .io_cfg_addr(pes_0_io_cfg_addr),
    .io_cfg_data(pes_0_io_cfg_data),
    .io_en(pes_0_io_en),
    .io_in_0(pes_0_io_in_0),
    .io_in_1(pes_0_io_in_1),
    .io_in_2(pes_0_io_in_2),
    .io_in_3(pes_0_io_in_3),
    .io_in_4(pes_0_io_in_4),
    .io_in_5(pes_0_io_in_5),
    .io_in_6(pes_0_io_in_6),
    .io_in_7(pes_0_io_in_7),
    .io_out_0(pes_0_io_out_0)
  );
  GPE_1 pes_1 ( // @[CGRA.scala 242:20]
    .clock(pes_1_clock),
    .reset(pes_1_reset),
    .io_cfg_en(pes_1_io_cfg_en),
    .io_cfg_addr(pes_1_io_cfg_addr),
    .io_cfg_data(pes_1_io_cfg_data),
    .io_en(pes_1_io_en),
    .io_in_0(pes_1_io_in_0),
    .io_in_1(pes_1_io_in_1),
    .io_in_2(pes_1_io_in_2),
    .io_in_3(pes_1_io_in_3),
    .io_in_4(pes_1_io_in_4),
    .io_in_5(pes_1_io_in_5),
    .io_in_6(pes_1_io_in_6),
    .io_in_7(pes_1_io_in_7),
    .io_out_0(pes_1_io_out_0)
  );
  GPE_2 pes_2 ( // @[CGRA.scala 242:20]
    .clock(pes_2_clock),
    .reset(pes_2_reset),
    .io_cfg_en(pes_2_io_cfg_en),
    .io_cfg_addr(pes_2_io_cfg_addr),
    .io_cfg_data(pes_2_io_cfg_data),
    .io_en(pes_2_io_en),
    .io_in_0(pes_2_io_in_0),
    .io_in_1(pes_2_io_in_1),
    .io_in_2(pes_2_io_in_2),
    .io_in_3(pes_2_io_in_3),
    .io_in_4(pes_2_io_in_4),
    .io_in_5(pes_2_io_in_5),
    .io_in_6(pes_2_io_in_6),
    .io_in_7(pes_2_io_in_7),
    .io_out_0(pes_2_io_out_0)
  );
  GPE_3 pes_3 ( // @[CGRA.scala 242:20]
    .clock(pes_3_clock),
    .reset(pes_3_reset),
    .io_cfg_en(pes_3_io_cfg_en),
    .io_cfg_addr(pes_3_io_cfg_addr),
    .io_cfg_data(pes_3_io_cfg_data),
    .io_en(pes_3_io_en),
    .io_in_0(pes_3_io_in_0),
    .io_in_1(pes_3_io_in_1),
    .io_in_2(pes_3_io_in_2),
    .io_in_3(pes_3_io_in_3),
    .io_in_4(pes_3_io_in_4),
    .io_in_5(pes_3_io_in_5),
    .io_in_6(pes_3_io_in_6),
    .io_in_7(pes_3_io_in_7),
    .io_out_0(pes_3_io_out_0)
  );
  GPE_4 pes_4 ( // @[CGRA.scala 242:20]
    .clock(pes_4_clock),
    .reset(pes_4_reset),
    .io_cfg_en(pes_4_io_cfg_en),
    .io_cfg_addr(pes_4_io_cfg_addr),
    .io_cfg_data(pes_4_io_cfg_data),
    .io_en(pes_4_io_en),
    .io_in_0(pes_4_io_in_0),
    .io_in_1(pes_4_io_in_1),
    .io_in_2(pes_4_io_in_2),
    .io_in_3(pes_4_io_in_3),
    .io_in_4(pes_4_io_in_4),
    .io_in_5(pes_4_io_in_5),
    .io_in_6(pes_4_io_in_6),
    .io_in_7(pes_4_io_in_7),
    .io_out_0(pes_4_io_out_0)
  );
  GPE_5 pes_5 ( // @[CGRA.scala 242:20]
    .clock(pes_5_clock),
    .reset(pes_5_reset),
    .io_cfg_en(pes_5_io_cfg_en),
    .io_cfg_addr(pes_5_io_cfg_addr),
    .io_cfg_data(pes_5_io_cfg_data),
    .io_en(pes_5_io_en),
    .io_in_0(pes_5_io_in_0),
    .io_in_1(pes_5_io_in_1),
    .io_in_2(pes_5_io_in_2),
    .io_in_3(pes_5_io_in_3),
    .io_in_4(pes_5_io_in_4),
    .io_in_5(pes_5_io_in_5),
    .io_in_6(pes_5_io_in_6),
    .io_in_7(pes_5_io_in_7),
    .io_out_0(pes_5_io_out_0)
  );
  GPE_6 pes_6 ( // @[CGRA.scala 242:20]
    .clock(pes_6_clock),
    .reset(pes_6_reset),
    .io_cfg_en(pes_6_io_cfg_en),
    .io_cfg_addr(pes_6_io_cfg_addr),
    .io_cfg_data(pes_6_io_cfg_data),
    .io_en(pes_6_io_en),
    .io_in_0(pes_6_io_in_0),
    .io_in_1(pes_6_io_in_1),
    .io_in_2(pes_6_io_in_2),
    .io_in_3(pes_6_io_in_3),
    .io_in_4(pes_6_io_in_4),
    .io_in_5(pes_6_io_in_5),
    .io_in_6(pes_6_io_in_6),
    .io_in_7(pes_6_io_in_7),
    .io_out_0(pes_6_io_out_0)
  );
  GPE_7 pes_7 ( // @[CGRA.scala 242:20]
    .clock(pes_7_clock),
    .reset(pes_7_reset),
    .io_cfg_en(pes_7_io_cfg_en),
    .io_cfg_addr(pes_7_io_cfg_addr),
    .io_cfg_data(pes_7_io_cfg_data),
    .io_en(pes_7_io_en),
    .io_in_0(pes_7_io_in_0),
    .io_in_1(pes_7_io_in_1),
    .io_in_2(pes_7_io_in_2),
    .io_in_3(pes_7_io_in_3),
    .io_in_4(pes_7_io_in_4),
    .io_in_5(pes_7_io_in_5),
    .io_in_6(pes_7_io_in_6),
    .io_in_7(pes_7_io_in_7),
    .io_out_0(pes_7_io_out_0)
  );
  GPE_8 pes_8 ( // @[CGRA.scala 242:20]
    .clock(pes_8_clock),
    .reset(pes_8_reset),
    .io_cfg_en(pes_8_io_cfg_en),
    .io_cfg_addr(pes_8_io_cfg_addr),
    .io_cfg_data(pes_8_io_cfg_data),
    .io_en(pes_8_io_en),
    .io_in_0(pes_8_io_in_0),
    .io_in_1(pes_8_io_in_1),
    .io_in_2(pes_8_io_in_2),
    .io_in_3(pes_8_io_in_3),
    .io_in_4(pes_8_io_in_4),
    .io_in_5(pes_8_io_in_5),
    .io_in_6(pes_8_io_in_6),
    .io_in_7(pes_8_io_in_7),
    .io_out_0(pes_8_io_out_0)
  );
  GPE_9 pes_9 ( // @[CGRA.scala 242:20]
    .clock(pes_9_clock),
    .reset(pes_9_reset),
    .io_cfg_en(pes_9_io_cfg_en),
    .io_cfg_addr(pes_9_io_cfg_addr),
    .io_cfg_data(pes_9_io_cfg_data),
    .io_en(pes_9_io_en),
    .io_in_0(pes_9_io_in_0),
    .io_in_1(pes_9_io_in_1),
    .io_in_2(pes_9_io_in_2),
    .io_in_3(pes_9_io_in_3),
    .io_in_4(pes_9_io_in_4),
    .io_in_5(pes_9_io_in_5),
    .io_in_6(pes_9_io_in_6),
    .io_in_7(pes_9_io_in_7),
    .io_out_0(pes_9_io_out_0)
  );
  GPE_10 pes_10 ( // @[CGRA.scala 242:20]
    .clock(pes_10_clock),
    .reset(pes_10_reset),
    .io_cfg_en(pes_10_io_cfg_en),
    .io_cfg_addr(pes_10_io_cfg_addr),
    .io_cfg_data(pes_10_io_cfg_data),
    .io_en(pes_10_io_en),
    .io_in_0(pes_10_io_in_0),
    .io_in_1(pes_10_io_in_1),
    .io_in_2(pes_10_io_in_2),
    .io_in_3(pes_10_io_in_3),
    .io_in_4(pes_10_io_in_4),
    .io_in_5(pes_10_io_in_5),
    .io_in_6(pes_10_io_in_6),
    .io_in_7(pes_10_io_in_7),
    .io_out_0(pes_10_io_out_0)
  );
  GPE_11 pes_11 ( // @[CGRA.scala 242:20]
    .clock(pes_11_clock),
    .reset(pes_11_reset),
    .io_cfg_en(pes_11_io_cfg_en),
    .io_cfg_addr(pes_11_io_cfg_addr),
    .io_cfg_data(pes_11_io_cfg_data),
    .io_en(pes_11_io_en),
    .io_in_0(pes_11_io_in_0),
    .io_in_1(pes_11_io_in_1),
    .io_in_2(pes_11_io_in_2),
    .io_in_3(pes_11_io_in_3),
    .io_in_4(pes_11_io_in_4),
    .io_in_5(pes_11_io_in_5),
    .io_in_6(pes_11_io_in_6),
    .io_in_7(pes_11_io_in_7),
    .io_out_0(pes_11_io_out_0)
  );
  GPE_12 pes_12 ( // @[CGRA.scala 242:20]
    .clock(pes_12_clock),
    .reset(pes_12_reset),
    .io_cfg_en(pes_12_io_cfg_en),
    .io_cfg_addr(pes_12_io_cfg_addr),
    .io_cfg_data(pes_12_io_cfg_data),
    .io_en(pes_12_io_en),
    .io_in_0(pes_12_io_in_0),
    .io_in_1(pes_12_io_in_1),
    .io_in_2(pes_12_io_in_2),
    .io_in_3(pes_12_io_in_3),
    .io_in_4(pes_12_io_in_4),
    .io_in_5(pes_12_io_in_5),
    .io_in_6(pes_12_io_in_6),
    .io_in_7(pes_12_io_in_7),
    .io_out_0(pes_12_io_out_0)
  );
  GPE_13 pes_13 ( // @[CGRA.scala 242:20]
    .clock(pes_13_clock),
    .reset(pes_13_reset),
    .io_cfg_en(pes_13_io_cfg_en),
    .io_cfg_addr(pes_13_io_cfg_addr),
    .io_cfg_data(pes_13_io_cfg_data),
    .io_en(pes_13_io_en),
    .io_in_0(pes_13_io_in_0),
    .io_in_1(pes_13_io_in_1),
    .io_in_2(pes_13_io_in_2),
    .io_in_3(pes_13_io_in_3),
    .io_in_4(pes_13_io_in_4),
    .io_in_5(pes_13_io_in_5),
    .io_in_6(pes_13_io_in_6),
    .io_in_7(pes_13_io_in_7),
    .io_out_0(pes_13_io_out_0)
  );
  GPE_14 pes_14 ( // @[CGRA.scala 242:20]
    .clock(pes_14_clock),
    .reset(pes_14_reset),
    .io_cfg_en(pes_14_io_cfg_en),
    .io_cfg_addr(pes_14_io_cfg_addr),
    .io_cfg_data(pes_14_io_cfg_data),
    .io_en(pes_14_io_en),
    .io_in_0(pes_14_io_in_0),
    .io_in_1(pes_14_io_in_1),
    .io_in_2(pes_14_io_in_2),
    .io_in_3(pes_14_io_in_3),
    .io_in_4(pes_14_io_in_4),
    .io_in_5(pes_14_io_in_5),
    .io_in_6(pes_14_io_in_6),
    .io_in_7(pes_14_io_in_7),
    .io_out_0(pes_14_io_out_0)
  );
  GPE_15 pes_15 ( // @[CGRA.scala 242:20]
    .clock(pes_15_clock),
    .reset(pes_15_reset),
    .io_cfg_en(pes_15_io_cfg_en),
    .io_cfg_addr(pes_15_io_cfg_addr),
    .io_cfg_data(pes_15_io_cfg_data),
    .io_en(pes_15_io_en),
    .io_in_0(pes_15_io_in_0),
    .io_in_1(pes_15_io_in_1),
    .io_in_2(pes_15_io_in_2),
    .io_in_3(pes_15_io_in_3),
    .io_in_4(pes_15_io_in_4),
    .io_in_5(pes_15_io_in_5),
    .io_in_6(pes_15_io_in_6),
    .io_in_7(pes_15_io_in_7),
    .io_out_0(pes_15_io_out_0)
  );
  GPE_16 pes_16 ( // @[CGRA.scala 242:20]
    .clock(pes_16_clock),
    .reset(pes_16_reset),
    .io_cfg_en(pes_16_io_cfg_en),
    .io_cfg_addr(pes_16_io_cfg_addr),
    .io_cfg_data(pes_16_io_cfg_data),
    .io_en(pes_16_io_en),
    .io_in_0(pes_16_io_in_0),
    .io_in_1(pes_16_io_in_1),
    .io_in_2(pes_16_io_in_2),
    .io_in_3(pes_16_io_in_3),
    .io_in_4(pes_16_io_in_4),
    .io_in_5(pes_16_io_in_5),
    .io_in_6(pes_16_io_in_6),
    .io_in_7(pes_16_io_in_7),
    .io_out_0(pes_16_io_out_0)
  );
  GPE_17 pes_17 ( // @[CGRA.scala 242:20]
    .clock(pes_17_clock),
    .reset(pes_17_reset),
    .io_cfg_en(pes_17_io_cfg_en),
    .io_cfg_addr(pes_17_io_cfg_addr),
    .io_cfg_data(pes_17_io_cfg_data),
    .io_en(pes_17_io_en),
    .io_in_0(pes_17_io_in_0),
    .io_in_1(pes_17_io_in_1),
    .io_in_2(pes_17_io_in_2),
    .io_in_3(pes_17_io_in_3),
    .io_in_4(pes_17_io_in_4),
    .io_in_5(pes_17_io_in_5),
    .io_in_6(pes_17_io_in_6),
    .io_in_7(pes_17_io_in_7),
    .io_out_0(pes_17_io_out_0)
  );
  GPE_18 pes_18 ( // @[CGRA.scala 242:20]
    .clock(pes_18_clock),
    .reset(pes_18_reset),
    .io_cfg_en(pes_18_io_cfg_en),
    .io_cfg_addr(pes_18_io_cfg_addr),
    .io_cfg_data(pes_18_io_cfg_data),
    .io_en(pes_18_io_en),
    .io_in_0(pes_18_io_in_0),
    .io_in_1(pes_18_io_in_1),
    .io_in_2(pes_18_io_in_2),
    .io_in_3(pes_18_io_in_3),
    .io_in_4(pes_18_io_in_4),
    .io_in_5(pes_18_io_in_5),
    .io_in_6(pes_18_io_in_6),
    .io_in_7(pes_18_io_in_7),
    .io_out_0(pes_18_io_out_0)
  );
  GPE_19 pes_19 ( // @[CGRA.scala 242:20]
    .clock(pes_19_clock),
    .reset(pes_19_reset),
    .io_cfg_en(pes_19_io_cfg_en),
    .io_cfg_addr(pes_19_io_cfg_addr),
    .io_cfg_data(pes_19_io_cfg_data),
    .io_en(pes_19_io_en),
    .io_in_0(pes_19_io_in_0),
    .io_in_1(pes_19_io_in_1),
    .io_in_2(pes_19_io_in_2),
    .io_in_3(pes_19_io_in_3),
    .io_in_4(pes_19_io_in_4),
    .io_in_5(pes_19_io_in_5),
    .io_in_6(pes_19_io_in_6),
    .io_in_7(pes_19_io_in_7),
    .io_out_0(pes_19_io_out_0)
  );
  GPE_20 pes_20 ( // @[CGRA.scala 242:20]
    .clock(pes_20_clock),
    .reset(pes_20_reset),
    .io_cfg_en(pes_20_io_cfg_en),
    .io_cfg_addr(pes_20_io_cfg_addr),
    .io_cfg_data(pes_20_io_cfg_data),
    .io_en(pes_20_io_en),
    .io_in_0(pes_20_io_in_0),
    .io_in_1(pes_20_io_in_1),
    .io_in_2(pes_20_io_in_2),
    .io_in_3(pes_20_io_in_3),
    .io_in_4(pes_20_io_in_4),
    .io_in_5(pes_20_io_in_5),
    .io_in_6(pes_20_io_in_6),
    .io_in_7(pes_20_io_in_7),
    .io_out_0(pes_20_io_out_0)
  );
  GPE_21 pes_21 ( // @[CGRA.scala 242:20]
    .clock(pes_21_clock),
    .reset(pes_21_reset),
    .io_cfg_en(pes_21_io_cfg_en),
    .io_cfg_addr(pes_21_io_cfg_addr),
    .io_cfg_data(pes_21_io_cfg_data),
    .io_en(pes_21_io_en),
    .io_in_0(pes_21_io_in_0),
    .io_in_1(pes_21_io_in_1),
    .io_in_2(pes_21_io_in_2),
    .io_in_3(pes_21_io_in_3),
    .io_in_4(pes_21_io_in_4),
    .io_in_5(pes_21_io_in_5),
    .io_in_6(pes_21_io_in_6),
    .io_in_7(pes_21_io_in_7),
    .io_out_0(pes_21_io_out_0)
  );
  GPE_22 pes_22 ( // @[CGRA.scala 242:20]
    .clock(pes_22_clock),
    .reset(pes_22_reset),
    .io_cfg_en(pes_22_io_cfg_en),
    .io_cfg_addr(pes_22_io_cfg_addr),
    .io_cfg_data(pes_22_io_cfg_data),
    .io_en(pes_22_io_en),
    .io_in_0(pes_22_io_in_0),
    .io_in_1(pes_22_io_in_1),
    .io_in_2(pes_22_io_in_2),
    .io_in_3(pes_22_io_in_3),
    .io_in_4(pes_22_io_in_4),
    .io_in_5(pes_22_io_in_5),
    .io_in_6(pes_22_io_in_6),
    .io_in_7(pes_22_io_in_7),
    .io_out_0(pes_22_io_out_0)
  );
  GPE_23 pes_23 ( // @[CGRA.scala 242:20]
    .clock(pes_23_clock),
    .reset(pes_23_reset),
    .io_cfg_en(pes_23_io_cfg_en),
    .io_cfg_addr(pes_23_io_cfg_addr),
    .io_cfg_data(pes_23_io_cfg_data),
    .io_en(pes_23_io_en),
    .io_in_0(pes_23_io_in_0),
    .io_in_1(pes_23_io_in_1),
    .io_in_2(pes_23_io_in_2),
    .io_in_3(pes_23_io_in_3),
    .io_in_4(pes_23_io_in_4),
    .io_in_5(pes_23_io_in_5),
    .io_in_6(pes_23_io_in_6),
    .io_in_7(pes_23_io_in_7),
    .io_out_0(pes_23_io_out_0)
  );
  GPE_24 pes_24 ( // @[CGRA.scala 242:20]
    .clock(pes_24_clock),
    .reset(pes_24_reset),
    .io_cfg_en(pes_24_io_cfg_en),
    .io_cfg_addr(pes_24_io_cfg_addr),
    .io_cfg_data(pes_24_io_cfg_data),
    .io_en(pes_24_io_en),
    .io_in_0(pes_24_io_in_0),
    .io_in_1(pes_24_io_in_1),
    .io_in_2(pes_24_io_in_2),
    .io_in_3(pes_24_io_in_3),
    .io_in_4(pes_24_io_in_4),
    .io_in_5(pes_24_io_in_5),
    .io_in_6(pes_24_io_in_6),
    .io_in_7(pes_24_io_in_7),
    .io_out_0(pes_24_io_out_0)
  );
  GPE_25 pes_25 ( // @[CGRA.scala 242:20]
    .clock(pes_25_clock),
    .reset(pes_25_reset),
    .io_cfg_en(pes_25_io_cfg_en),
    .io_cfg_addr(pes_25_io_cfg_addr),
    .io_cfg_data(pes_25_io_cfg_data),
    .io_en(pes_25_io_en),
    .io_in_0(pes_25_io_in_0),
    .io_in_1(pes_25_io_in_1),
    .io_in_2(pes_25_io_in_2),
    .io_in_3(pes_25_io_in_3),
    .io_in_4(pes_25_io_in_4),
    .io_in_5(pes_25_io_in_5),
    .io_in_6(pes_25_io_in_6),
    .io_in_7(pes_25_io_in_7),
    .io_out_0(pes_25_io_out_0)
  );
  GPE_26 pes_26 ( // @[CGRA.scala 242:20]
    .clock(pes_26_clock),
    .reset(pes_26_reset),
    .io_cfg_en(pes_26_io_cfg_en),
    .io_cfg_addr(pes_26_io_cfg_addr),
    .io_cfg_data(pes_26_io_cfg_data),
    .io_en(pes_26_io_en),
    .io_in_0(pes_26_io_in_0),
    .io_in_1(pes_26_io_in_1),
    .io_in_2(pes_26_io_in_2),
    .io_in_3(pes_26_io_in_3),
    .io_in_4(pes_26_io_in_4),
    .io_in_5(pes_26_io_in_5),
    .io_in_6(pes_26_io_in_6),
    .io_in_7(pes_26_io_in_7),
    .io_out_0(pes_26_io_out_0)
  );
  GPE_27 pes_27 ( // @[CGRA.scala 242:20]
    .clock(pes_27_clock),
    .reset(pes_27_reset),
    .io_cfg_en(pes_27_io_cfg_en),
    .io_cfg_addr(pes_27_io_cfg_addr),
    .io_cfg_data(pes_27_io_cfg_data),
    .io_en(pes_27_io_en),
    .io_in_0(pes_27_io_in_0),
    .io_in_1(pes_27_io_in_1),
    .io_in_2(pes_27_io_in_2),
    .io_in_3(pes_27_io_in_3),
    .io_in_4(pes_27_io_in_4),
    .io_in_5(pes_27_io_in_5),
    .io_in_6(pes_27_io_in_6),
    .io_in_7(pes_27_io_in_7),
    .io_out_0(pes_27_io_out_0)
  );
  GPE_28 pes_28 ( // @[CGRA.scala 242:20]
    .clock(pes_28_clock),
    .reset(pes_28_reset),
    .io_cfg_en(pes_28_io_cfg_en),
    .io_cfg_addr(pes_28_io_cfg_addr),
    .io_cfg_data(pes_28_io_cfg_data),
    .io_en(pes_28_io_en),
    .io_in_0(pes_28_io_in_0),
    .io_in_1(pes_28_io_in_1),
    .io_in_2(pes_28_io_in_2),
    .io_in_3(pes_28_io_in_3),
    .io_in_4(pes_28_io_in_4),
    .io_in_5(pes_28_io_in_5),
    .io_in_6(pes_28_io_in_6),
    .io_in_7(pes_28_io_in_7),
    .io_out_0(pes_28_io_out_0)
  );
  GPE_29 pes_29 ( // @[CGRA.scala 242:20]
    .clock(pes_29_clock),
    .reset(pes_29_reset),
    .io_cfg_en(pes_29_io_cfg_en),
    .io_cfg_addr(pes_29_io_cfg_addr),
    .io_cfg_data(pes_29_io_cfg_data),
    .io_en(pes_29_io_en),
    .io_in_0(pes_29_io_in_0),
    .io_in_1(pes_29_io_in_1),
    .io_in_2(pes_29_io_in_2),
    .io_in_3(pes_29_io_in_3),
    .io_in_4(pes_29_io_in_4),
    .io_in_5(pes_29_io_in_5),
    .io_in_6(pes_29_io_in_6),
    .io_in_7(pes_29_io_in_7),
    .io_out_0(pes_29_io_out_0)
  );
  GPE_30 pes_30 ( // @[CGRA.scala 242:20]
    .clock(pes_30_clock),
    .reset(pes_30_reset),
    .io_cfg_en(pes_30_io_cfg_en),
    .io_cfg_addr(pes_30_io_cfg_addr),
    .io_cfg_data(pes_30_io_cfg_data),
    .io_en(pes_30_io_en),
    .io_in_0(pes_30_io_in_0),
    .io_in_1(pes_30_io_in_1),
    .io_in_2(pes_30_io_in_2),
    .io_in_3(pes_30_io_in_3),
    .io_in_4(pes_30_io_in_4),
    .io_in_5(pes_30_io_in_5),
    .io_in_6(pes_30_io_in_6),
    .io_in_7(pes_30_io_in_7),
    .io_out_0(pes_30_io_out_0)
  );
  GPE_31 pes_31 ( // @[CGRA.scala 242:20]
    .clock(pes_31_clock),
    .reset(pes_31_reset),
    .io_cfg_en(pes_31_io_cfg_en),
    .io_cfg_addr(pes_31_io_cfg_addr),
    .io_cfg_data(pes_31_io_cfg_data),
    .io_en(pes_31_io_en),
    .io_in_0(pes_31_io_in_0),
    .io_in_1(pes_31_io_in_1),
    .io_in_2(pes_31_io_in_2),
    .io_in_3(pes_31_io_in_3),
    .io_in_4(pes_31_io_in_4),
    .io_in_5(pes_31_io_in_5),
    .io_in_6(pes_31_io_in_6),
    .io_in_7(pes_31_io_in_7),
    .io_out_0(pes_31_io_out_0)
  );
  GPE_32 pes_32 ( // @[CGRA.scala 242:20]
    .clock(pes_32_clock),
    .reset(pes_32_reset),
    .io_cfg_en(pes_32_io_cfg_en),
    .io_cfg_addr(pes_32_io_cfg_addr),
    .io_cfg_data(pes_32_io_cfg_data),
    .io_en(pes_32_io_en),
    .io_in_0(pes_32_io_in_0),
    .io_in_1(pes_32_io_in_1),
    .io_in_2(pes_32_io_in_2),
    .io_in_3(pes_32_io_in_3),
    .io_in_4(pes_32_io_in_4),
    .io_in_5(pes_32_io_in_5),
    .io_in_6(pes_32_io_in_6),
    .io_in_7(pes_32_io_in_7),
    .io_out_0(pes_32_io_out_0)
  );
  GPE_33 pes_33 ( // @[CGRA.scala 242:20]
    .clock(pes_33_clock),
    .reset(pes_33_reset),
    .io_cfg_en(pes_33_io_cfg_en),
    .io_cfg_addr(pes_33_io_cfg_addr),
    .io_cfg_data(pes_33_io_cfg_data),
    .io_en(pes_33_io_en),
    .io_in_0(pes_33_io_in_0),
    .io_in_1(pes_33_io_in_1),
    .io_in_2(pes_33_io_in_2),
    .io_in_3(pes_33_io_in_3),
    .io_in_4(pes_33_io_in_4),
    .io_in_5(pes_33_io_in_5),
    .io_in_6(pes_33_io_in_6),
    .io_in_7(pes_33_io_in_7),
    .io_out_0(pes_33_io_out_0)
  );
  GPE_34 pes_34 ( // @[CGRA.scala 242:20]
    .clock(pes_34_clock),
    .reset(pes_34_reset),
    .io_cfg_en(pes_34_io_cfg_en),
    .io_cfg_addr(pes_34_io_cfg_addr),
    .io_cfg_data(pes_34_io_cfg_data),
    .io_en(pes_34_io_en),
    .io_in_0(pes_34_io_in_0),
    .io_in_1(pes_34_io_in_1),
    .io_in_2(pes_34_io_in_2),
    .io_in_3(pes_34_io_in_3),
    .io_in_4(pes_34_io_in_4),
    .io_in_5(pes_34_io_in_5),
    .io_in_6(pes_34_io_in_6),
    .io_in_7(pes_34_io_in_7),
    .io_out_0(pes_34_io_out_0)
  );
  GPE_35 pes_35 ( // @[CGRA.scala 242:20]
    .clock(pes_35_clock),
    .reset(pes_35_reset),
    .io_cfg_en(pes_35_io_cfg_en),
    .io_cfg_addr(pes_35_io_cfg_addr),
    .io_cfg_data(pes_35_io_cfg_data),
    .io_en(pes_35_io_en),
    .io_in_0(pes_35_io_in_0),
    .io_in_1(pes_35_io_in_1),
    .io_in_2(pes_35_io_in_2),
    .io_in_3(pes_35_io_in_3),
    .io_in_4(pes_35_io_in_4),
    .io_in_5(pes_35_io_in_5),
    .io_in_6(pes_35_io_in_6),
    .io_in_7(pes_35_io_in_7),
    .io_out_0(pes_35_io_out_0)
  );
  GPE_36 pes_36 ( // @[CGRA.scala 242:20]
    .clock(pes_36_clock),
    .reset(pes_36_reset),
    .io_cfg_en(pes_36_io_cfg_en),
    .io_cfg_addr(pes_36_io_cfg_addr),
    .io_cfg_data(pes_36_io_cfg_data),
    .io_en(pes_36_io_en),
    .io_in_0(pes_36_io_in_0),
    .io_in_1(pes_36_io_in_1),
    .io_in_2(pes_36_io_in_2),
    .io_in_3(pes_36_io_in_3),
    .io_in_4(pes_36_io_in_4),
    .io_in_5(pes_36_io_in_5),
    .io_in_6(pes_36_io_in_6),
    .io_in_7(pes_36_io_in_7),
    .io_out_0(pes_36_io_out_0)
  );
  GPE_37 pes_37 ( // @[CGRA.scala 242:20]
    .clock(pes_37_clock),
    .reset(pes_37_reset),
    .io_cfg_en(pes_37_io_cfg_en),
    .io_cfg_addr(pes_37_io_cfg_addr),
    .io_cfg_data(pes_37_io_cfg_data),
    .io_en(pes_37_io_en),
    .io_in_0(pes_37_io_in_0),
    .io_in_1(pes_37_io_in_1),
    .io_in_2(pes_37_io_in_2),
    .io_in_3(pes_37_io_in_3),
    .io_in_4(pes_37_io_in_4),
    .io_in_5(pes_37_io_in_5),
    .io_in_6(pes_37_io_in_6),
    .io_in_7(pes_37_io_in_7),
    .io_out_0(pes_37_io_out_0)
  );
  GPE_38 pes_38 ( // @[CGRA.scala 242:20]
    .clock(pes_38_clock),
    .reset(pes_38_reset),
    .io_cfg_en(pes_38_io_cfg_en),
    .io_cfg_addr(pes_38_io_cfg_addr),
    .io_cfg_data(pes_38_io_cfg_data),
    .io_en(pes_38_io_en),
    .io_in_0(pes_38_io_in_0),
    .io_in_1(pes_38_io_in_1),
    .io_in_2(pes_38_io_in_2),
    .io_in_3(pes_38_io_in_3),
    .io_in_4(pes_38_io_in_4),
    .io_in_5(pes_38_io_in_5),
    .io_in_6(pes_38_io_in_6),
    .io_in_7(pes_38_io_in_7),
    .io_out_0(pes_38_io_out_0)
  );
  GPE_39 pes_39 ( // @[CGRA.scala 242:20]
    .clock(pes_39_clock),
    .reset(pes_39_reset),
    .io_cfg_en(pes_39_io_cfg_en),
    .io_cfg_addr(pes_39_io_cfg_addr),
    .io_cfg_data(pes_39_io_cfg_data),
    .io_en(pes_39_io_en),
    .io_in_0(pes_39_io_in_0),
    .io_in_1(pes_39_io_in_1),
    .io_in_2(pes_39_io_in_2),
    .io_in_3(pes_39_io_in_3),
    .io_in_4(pes_39_io_in_4),
    .io_in_5(pes_39_io_in_5),
    .io_in_6(pes_39_io_in_6),
    .io_in_7(pes_39_io_in_7),
    .io_out_0(pes_39_io_out_0)
  );
  GPE_40 pes_40 ( // @[CGRA.scala 242:20]
    .clock(pes_40_clock),
    .reset(pes_40_reset),
    .io_cfg_en(pes_40_io_cfg_en),
    .io_cfg_addr(pes_40_io_cfg_addr),
    .io_cfg_data(pes_40_io_cfg_data),
    .io_en(pes_40_io_en),
    .io_in_0(pes_40_io_in_0),
    .io_in_1(pes_40_io_in_1),
    .io_in_2(pes_40_io_in_2),
    .io_in_3(pes_40_io_in_3),
    .io_in_4(pes_40_io_in_4),
    .io_in_5(pes_40_io_in_5),
    .io_in_6(pes_40_io_in_6),
    .io_in_7(pes_40_io_in_7),
    .io_out_0(pes_40_io_out_0)
  );
  GPE_41 pes_41 ( // @[CGRA.scala 242:20]
    .clock(pes_41_clock),
    .reset(pes_41_reset),
    .io_cfg_en(pes_41_io_cfg_en),
    .io_cfg_addr(pes_41_io_cfg_addr),
    .io_cfg_data(pes_41_io_cfg_data),
    .io_en(pes_41_io_en),
    .io_in_0(pes_41_io_in_0),
    .io_in_1(pes_41_io_in_1),
    .io_in_2(pes_41_io_in_2),
    .io_in_3(pes_41_io_in_3),
    .io_in_4(pes_41_io_in_4),
    .io_in_5(pes_41_io_in_5),
    .io_in_6(pes_41_io_in_6),
    .io_in_7(pes_41_io_in_7),
    .io_out_0(pes_41_io_out_0)
  );
  GPE_42 pes_42 ( // @[CGRA.scala 242:20]
    .clock(pes_42_clock),
    .reset(pes_42_reset),
    .io_cfg_en(pes_42_io_cfg_en),
    .io_cfg_addr(pes_42_io_cfg_addr),
    .io_cfg_data(pes_42_io_cfg_data),
    .io_en(pes_42_io_en),
    .io_in_0(pes_42_io_in_0),
    .io_in_1(pes_42_io_in_1),
    .io_in_2(pes_42_io_in_2),
    .io_in_3(pes_42_io_in_3),
    .io_in_4(pes_42_io_in_4),
    .io_in_5(pes_42_io_in_5),
    .io_in_6(pes_42_io_in_6),
    .io_in_7(pes_42_io_in_7),
    .io_out_0(pes_42_io_out_0)
  );
  GPE_43 pes_43 ( // @[CGRA.scala 242:20]
    .clock(pes_43_clock),
    .reset(pes_43_reset),
    .io_cfg_en(pes_43_io_cfg_en),
    .io_cfg_addr(pes_43_io_cfg_addr),
    .io_cfg_data(pes_43_io_cfg_data),
    .io_en(pes_43_io_en),
    .io_in_0(pes_43_io_in_0),
    .io_in_1(pes_43_io_in_1),
    .io_in_2(pes_43_io_in_2),
    .io_in_3(pes_43_io_in_3),
    .io_in_4(pes_43_io_in_4),
    .io_in_5(pes_43_io_in_5),
    .io_in_6(pes_43_io_in_6),
    .io_in_7(pes_43_io_in_7),
    .io_out_0(pes_43_io_out_0)
  );
  GPE_44 pes_44 ( // @[CGRA.scala 242:20]
    .clock(pes_44_clock),
    .reset(pes_44_reset),
    .io_cfg_en(pes_44_io_cfg_en),
    .io_cfg_addr(pes_44_io_cfg_addr),
    .io_cfg_data(pes_44_io_cfg_data),
    .io_en(pes_44_io_en),
    .io_in_0(pes_44_io_in_0),
    .io_in_1(pes_44_io_in_1),
    .io_in_2(pes_44_io_in_2),
    .io_in_3(pes_44_io_in_3),
    .io_in_4(pes_44_io_in_4),
    .io_in_5(pes_44_io_in_5),
    .io_in_6(pes_44_io_in_6),
    .io_in_7(pes_44_io_in_7),
    .io_out_0(pes_44_io_out_0)
  );
  GPE_45 pes_45 ( // @[CGRA.scala 242:20]
    .clock(pes_45_clock),
    .reset(pes_45_reset),
    .io_cfg_en(pes_45_io_cfg_en),
    .io_cfg_addr(pes_45_io_cfg_addr),
    .io_cfg_data(pes_45_io_cfg_data),
    .io_en(pes_45_io_en),
    .io_in_0(pes_45_io_in_0),
    .io_in_1(pes_45_io_in_1),
    .io_in_2(pes_45_io_in_2),
    .io_in_3(pes_45_io_in_3),
    .io_in_4(pes_45_io_in_4),
    .io_in_5(pes_45_io_in_5),
    .io_in_6(pes_45_io_in_6),
    .io_in_7(pes_45_io_in_7),
    .io_out_0(pes_45_io_out_0)
  );
  GPE_46 pes_46 ( // @[CGRA.scala 242:20]
    .clock(pes_46_clock),
    .reset(pes_46_reset),
    .io_cfg_en(pes_46_io_cfg_en),
    .io_cfg_addr(pes_46_io_cfg_addr),
    .io_cfg_data(pes_46_io_cfg_data),
    .io_en(pes_46_io_en),
    .io_in_0(pes_46_io_in_0),
    .io_in_1(pes_46_io_in_1),
    .io_in_2(pes_46_io_in_2),
    .io_in_3(pes_46_io_in_3),
    .io_in_4(pes_46_io_in_4),
    .io_in_5(pes_46_io_in_5),
    .io_in_6(pes_46_io_in_6),
    .io_in_7(pes_46_io_in_7),
    .io_out_0(pes_46_io_out_0)
  );
  GPE_47 pes_47 ( // @[CGRA.scala 242:20]
    .clock(pes_47_clock),
    .reset(pes_47_reset),
    .io_cfg_en(pes_47_io_cfg_en),
    .io_cfg_addr(pes_47_io_cfg_addr),
    .io_cfg_data(pes_47_io_cfg_data),
    .io_en(pes_47_io_en),
    .io_in_0(pes_47_io_in_0),
    .io_in_1(pes_47_io_in_1),
    .io_in_2(pes_47_io_in_2),
    .io_in_3(pes_47_io_in_3),
    .io_in_4(pes_47_io_in_4),
    .io_in_5(pes_47_io_in_5),
    .io_in_6(pes_47_io_in_6),
    .io_in_7(pes_47_io_in_7),
    .io_out_0(pes_47_io_out_0)
  );
  GPE_48 pes_48 ( // @[CGRA.scala 242:20]
    .clock(pes_48_clock),
    .reset(pes_48_reset),
    .io_cfg_en(pes_48_io_cfg_en),
    .io_cfg_addr(pes_48_io_cfg_addr),
    .io_cfg_data(pes_48_io_cfg_data),
    .io_en(pes_48_io_en),
    .io_in_0(pes_48_io_in_0),
    .io_in_1(pes_48_io_in_1),
    .io_in_2(pes_48_io_in_2),
    .io_in_3(pes_48_io_in_3),
    .io_in_4(pes_48_io_in_4),
    .io_in_5(pes_48_io_in_5),
    .io_in_6(pes_48_io_in_6),
    .io_in_7(pes_48_io_in_7),
    .io_out_0(pes_48_io_out_0)
  );
  GPE_49 pes_49 ( // @[CGRA.scala 242:20]
    .clock(pes_49_clock),
    .reset(pes_49_reset),
    .io_cfg_en(pes_49_io_cfg_en),
    .io_cfg_addr(pes_49_io_cfg_addr),
    .io_cfg_data(pes_49_io_cfg_data),
    .io_en(pes_49_io_en),
    .io_in_0(pes_49_io_in_0),
    .io_in_1(pes_49_io_in_1),
    .io_in_2(pes_49_io_in_2),
    .io_in_3(pes_49_io_in_3),
    .io_in_4(pes_49_io_in_4),
    .io_in_5(pes_49_io_in_5),
    .io_in_6(pes_49_io_in_6),
    .io_in_7(pes_49_io_in_7),
    .io_out_0(pes_49_io_out_0)
  );
  GPE_50 pes_50 ( // @[CGRA.scala 242:20]
    .clock(pes_50_clock),
    .reset(pes_50_reset),
    .io_cfg_en(pes_50_io_cfg_en),
    .io_cfg_addr(pes_50_io_cfg_addr),
    .io_cfg_data(pes_50_io_cfg_data),
    .io_en(pes_50_io_en),
    .io_in_0(pes_50_io_in_0),
    .io_in_1(pes_50_io_in_1),
    .io_in_2(pes_50_io_in_2),
    .io_in_3(pes_50_io_in_3),
    .io_in_4(pes_50_io_in_4),
    .io_in_5(pes_50_io_in_5),
    .io_in_6(pes_50_io_in_6),
    .io_in_7(pes_50_io_in_7),
    .io_out_0(pes_50_io_out_0)
  );
  GPE_51 pes_51 ( // @[CGRA.scala 242:20]
    .clock(pes_51_clock),
    .reset(pes_51_reset),
    .io_cfg_en(pes_51_io_cfg_en),
    .io_cfg_addr(pes_51_io_cfg_addr),
    .io_cfg_data(pes_51_io_cfg_data),
    .io_en(pes_51_io_en),
    .io_in_0(pes_51_io_in_0),
    .io_in_1(pes_51_io_in_1),
    .io_in_2(pes_51_io_in_2),
    .io_in_3(pes_51_io_in_3),
    .io_in_4(pes_51_io_in_4),
    .io_in_5(pes_51_io_in_5),
    .io_in_6(pes_51_io_in_6),
    .io_in_7(pes_51_io_in_7),
    .io_out_0(pes_51_io_out_0)
  );
  GPE_52 pes_52 ( // @[CGRA.scala 242:20]
    .clock(pes_52_clock),
    .reset(pes_52_reset),
    .io_cfg_en(pes_52_io_cfg_en),
    .io_cfg_addr(pes_52_io_cfg_addr),
    .io_cfg_data(pes_52_io_cfg_data),
    .io_en(pes_52_io_en),
    .io_in_0(pes_52_io_in_0),
    .io_in_1(pes_52_io_in_1),
    .io_in_2(pes_52_io_in_2),
    .io_in_3(pes_52_io_in_3),
    .io_in_4(pes_52_io_in_4),
    .io_in_5(pes_52_io_in_5),
    .io_in_6(pes_52_io_in_6),
    .io_in_7(pes_52_io_in_7),
    .io_out_0(pes_52_io_out_0)
  );
  GPE_53 pes_53 ( // @[CGRA.scala 242:20]
    .clock(pes_53_clock),
    .reset(pes_53_reset),
    .io_cfg_en(pes_53_io_cfg_en),
    .io_cfg_addr(pes_53_io_cfg_addr),
    .io_cfg_data(pes_53_io_cfg_data),
    .io_en(pes_53_io_en),
    .io_in_0(pes_53_io_in_0),
    .io_in_1(pes_53_io_in_1),
    .io_in_2(pes_53_io_in_2),
    .io_in_3(pes_53_io_in_3),
    .io_in_4(pes_53_io_in_4),
    .io_in_5(pes_53_io_in_5),
    .io_in_6(pes_53_io_in_6),
    .io_in_7(pes_53_io_in_7),
    .io_out_0(pes_53_io_out_0)
  );
  GPE_54 pes_54 ( // @[CGRA.scala 242:20]
    .clock(pes_54_clock),
    .reset(pes_54_reset),
    .io_cfg_en(pes_54_io_cfg_en),
    .io_cfg_addr(pes_54_io_cfg_addr),
    .io_cfg_data(pes_54_io_cfg_data),
    .io_en(pes_54_io_en),
    .io_in_0(pes_54_io_in_0),
    .io_in_1(pes_54_io_in_1),
    .io_in_2(pes_54_io_in_2),
    .io_in_3(pes_54_io_in_3),
    .io_in_4(pes_54_io_in_4),
    .io_in_5(pes_54_io_in_5),
    .io_in_6(pes_54_io_in_6),
    .io_in_7(pes_54_io_in_7),
    .io_out_0(pes_54_io_out_0)
  );
  GPE_55 pes_55 ( // @[CGRA.scala 242:20]
    .clock(pes_55_clock),
    .reset(pes_55_reset),
    .io_cfg_en(pes_55_io_cfg_en),
    .io_cfg_addr(pes_55_io_cfg_addr),
    .io_cfg_data(pes_55_io_cfg_data),
    .io_en(pes_55_io_en),
    .io_in_0(pes_55_io_in_0),
    .io_in_1(pes_55_io_in_1),
    .io_in_2(pes_55_io_in_2),
    .io_in_3(pes_55_io_in_3),
    .io_in_4(pes_55_io_in_4),
    .io_in_5(pes_55_io_in_5),
    .io_in_6(pes_55_io_in_6),
    .io_in_7(pes_55_io_in_7),
    .io_out_0(pes_55_io_out_0)
  );
  GPE_56 pes_56 ( // @[CGRA.scala 242:20]
    .clock(pes_56_clock),
    .reset(pes_56_reset),
    .io_cfg_en(pes_56_io_cfg_en),
    .io_cfg_addr(pes_56_io_cfg_addr),
    .io_cfg_data(pes_56_io_cfg_data),
    .io_en(pes_56_io_en),
    .io_in_0(pes_56_io_in_0),
    .io_in_1(pes_56_io_in_1),
    .io_in_2(pes_56_io_in_2),
    .io_in_3(pes_56_io_in_3),
    .io_in_4(pes_56_io_in_4),
    .io_in_5(pes_56_io_in_5),
    .io_in_6(pes_56_io_in_6),
    .io_in_7(pes_56_io_in_7),
    .io_out_0(pes_56_io_out_0)
  );
  GIB gibs_0 ( // @[CGRA.scala 333:21]
    .clock(gibs_0_clock),
    .reset(gibs_0_reset),
    .io_cfg_en(gibs_0_io_cfg_en),
    .io_cfg_addr(gibs_0_io_cfg_addr),
    .io_cfg_data(gibs_0_io_cfg_data),
    .io_ipinNE_0(gibs_0_io_ipinNE_0),
    .io_opinNE_0(gibs_0_io_opinNE_0),
    .io_ipinSE_0(gibs_0_io_ipinSE_0),
    .io_ipinSE_1(gibs_0_io_ipinSE_1),
    .io_opinSE_0(gibs_0_io_opinSE_0),
    .io_ipinSW_0(gibs_0_io_ipinSW_0),
    .io_opinSW_0(gibs_0_io_opinSW_0),
    .io_itrackE_0(gibs_0_io_itrackE_0),
    .io_otrackE_0(gibs_0_io_otrackE_0),
    .io_itrackS_0(gibs_0_io_itrackS_0),
    .io_otrackS_0(gibs_0_io_otrackS_0)
  );
  GIB_1 gibs_1 ( // @[CGRA.scala 333:21]
    .clock(gibs_1_clock),
    .reset(gibs_1_reset),
    .io_cfg_en(gibs_1_io_cfg_en),
    .io_cfg_addr(gibs_1_io_cfg_addr),
    .io_cfg_data(gibs_1_io_cfg_data),
    .io_ipinNW_0(gibs_1_io_ipinNW_0),
    .io_opinNW_0(gibs_1_io_opinNW_0),
    .io_ipinNE_0(gibs_1_io_ipinNE_0),
    .io_opinNE_0(gibs_1_io_opinNE_0),
    .io_ipinSE_0(gibs_1_io_ipinSE_0),
    .io_ipinSE_1(gibs_1_io_ipinSE_1),
    .io_opinSE_0(gibs_1_io_opinSE_0),
    .io_ipinSW_0(gibs_1_io_ipinSW_0),
    .io_ipinSW_1(gibs_1_io_ipinSW_1),
    .io_opinSW_0(gibs_1_io_opinSW_0),
    .io_itrackW_0(gibs_1_io_itrackW_0),
    .io_otrackW_0(gibs_1_io_otrackW_0),
    .io_itrackE_0(gibs_1_io_itrackE_0),
    .io_otrackE_0(gibs_1_io_otrackE_0),
    .io_itrackS_0(gibs_1_io_itrackS_0),
    .io_otrackS_0(gibs_1_io_otrackS_0)
  );
  GIB_2 gibs_2 ( // @[CGRA.scala 333:21]
    .clock(gibs_2_clock),
    .reset(gibs_2_reset),
    .io_cfg_en(gibs_2_io_cfg_en),
    .io_cfg_addr(gibs_2_io_cfg_addr),
    .io_cfg_data(gibs_2_io_cfg_data),
    .io_ipinNW_0(gibs_2_io_ipinNW_0),
    .io_opinNW_0(gibs_2_io_opinNW_0),
    .io_ipinNE_0(gibs_2_io_ipinNE_0),
    .io_opinNE_0(gibs_2_io_opinNE_0),
    .io_ipinSE_0(gibs_2_io_ipinSE_0),
    .io_ipinSE_1(gibs_2_io_ipinSE_1),
    .io_opinSE_0(gibs_2_io_opinSE_0),
    .io_ipinSW_0(gibs_2_io_ipinSW_0),
    .io_ipinSW_1(gibs_2_io_ipinSW_1),
    .io_opinSW_0(gibs_2_io_opinSW_0),
    .io_itrackW_0(gibs_2_io_itrackW_0),
    .io_otrackW_0(gibs_2_io_otrackW_0),
    .io_itrackE_0(gibs_2_io_itrackE_0),
    .io_otrackE_0(gibs_2_io_otrackE_0),
    .io_itrackS_0(gibs_2_io_itrackS_0),
    .io_otrackS_0(gibs_2_io_otrackS_0)
  );
  GIB_3 gibs_3 ( // @[CGRA.scala 333:21]
    .clock(gibs_3_clock),
    .reset(gibs_3_reset),
    .io_cfg_en(gibs_3_io_cfg_en),
    .io_cfg_addr(gibs_3_io_cfg_addr),
    .io_cfg_data(gibs_3_io_cfg_data),
    .io_ipinNW_0(gibs_3_io_ipinNW_0),
    .io_opinNW_0(gibs_3_io_opinNW_0),
    .io_ipinSE_0(gibs_3_io_ipinSE_0),
    .io_opinSE_0(gibs_3_io_opinSE_0),
    .io_ipinSW_0(gibs_3_io_ipinSW_0),
    .io_ipinSW_1(gibs_3_io_ipinSW_1),
    .io_opinSW_0(gibs_3_io_opinSW_0),
    .io_itrackW_0(gibs_3_io_itrackW_0),
    .io_otrackW_0(gibs_3_io_otrackW_0),
    .io_itrackS_0(gibs_3_io_itrackS_0),
    .io_otrackS_0(gibs_3_io_otrackS_0)
  );
  GIB_4 gibs_4 ( // @[CGRA.scala 333:21]
    .clock(gibs_4_clock),
    .reset(gibs_4_reset),
    .io_cfg_en(gibs_4_io_cfg_en),
    .io_cfg_addr(gibs_4_io_cfg_addr),
    .io_cfg_data(gibs_4_io_cfg_data),
    .io_ipinNW_0(gibs_4_io_ipinNW_0),
    .io_opinNW_0(gibs_4_io_opinNW_0),
    .io_ipinNE_0(gibs_4_io_ipinNE_0),
    .io_ipinNE_1(gibs_4_io_ipinNE_1),
    .io_opinNE_0(gibs_4_io_opinNE_0),
    .io_ipinSE_0(gibs_4_io_ipinSE_0),
    .io_ipinSE_1(gibs_4_io_ipinSE_1),
    .io_opinSE_0(gibs_4_io_opinSE_0),
    .io_ipinSW_0(gibs_4_io_ipinSW_0),
    .io_opinSW_0(gibs_4_io_opinSW_0),
    .io_itrackN_0(gibs_4_io_itrackN_0),
    .io_otrackN_0(gibs_4_io_otrackN_0),
    .io_itrackE_0(gibs_4_io_itrackE_0),
    .io_otrackE_0(gibs_4_io_otrackE_0),
    .io_itrackS_0(gibs_4_io_itrackS_0),
    .io_otrackS_0(gibs_4_io_otrackS_0)
  );
  GIB_5 gibs_5 ( // @[CGRA.scala 333:21]
    .clock(gibs_5_clock),
    .reset(gibs_5_reset),
    .io_cfg_en(gibs_5_io_cfg_en),
    .io_cfg_addr(gibs_5_io_cfg_addr),
    .io_cfg_data(gibs_5_io_cfg_data),
    .io_ipinNW_0(gibs_5_io_ipinNW_0),
    .io_ipinNW_1(gibs_5_io_ipinNW_1),
    .io_opinNW_0(gibs_5_io_opinNW_0),
    .io_ipinNE_0(gibs_5_io_ipinNE_0),
    .io_ipinNE_1(gibs_5_io_ipinNE_1),
    .io_opinNE_0(gibs_5_io_opinNE_0),
    .io_ipinSE_0(gibs_5_io_ipinSE_0),
    .io_ipinSE_1(gibs_5_io_ipinSE_1),
    .io_opinSE_0(gibs_5_io_opinSE_0),
    .io_ipinSW_0(gibs_5_io_ipinSW_0),
    .io_ipinSW_1(gibs_5_io_ipinSW_1),
    .io_opinSW_0(gibs_5_io_opinSW_0),
    .io_itrackW_0(gibs_5_io_itrackW_0),
    .io_otrackW_0(gibs_5_io_otrackW_0),
    .io_itrackN_0(gibs_5_io_itrackN_0),
    .io_otrackN_0(gibs_5_io_otrackN_0),
    .io_itrackE_0(gibs_5_io_itrackE_0),
    .io_otrackE_0(gibs_5_io_otrackE_0),
    .io_itrackS_0(gibs_5_io_itrackS_0),
    .io_otrackS_0(gibs_5_io_otrackS_0)
  );
  GIB_6 gibs_6 ( // @[CGRA.scala 333:21]
    .clock(gibs_6_clock),
    .reset(gibs_6_reset),
    .io_cfg_en(gibs_6_io_cfg_en),
    .io_cfg_addr(gibs_6_io_cfg_addr),
    .io_cfg_data(gibs_6_io_cfg_data),
    .io_ipinNW_0(gibs_6_io_ipinNW_0),
    .io_ipinNW_1(gibs_6_io_ipinNW_1),
    .io_opinNW_0(gibs_6_io_opinNW_0),
    .io_ipinNE_0(gibs_6_io_ipinNE_0),
    .io_ipinNE_1(gibs_6_io_ipinNE_1),
    .io_opinNE_0(gibs_6_io_opinNE_0),
    .io_ipinSE_0(gibs_6_io_ipinSE_0),
    .io_ipinSE_1(gibs_6_io_ipinSE_1),
    .io_opinSE_0(gibs_6_io_opinSE_0),
    .io_ipinSW_0(gibs_6_io_ipinSW_0),
    .io_ipinSW_1(gibs_6_io_ipinSW_1),
    .io_opinSW_0(gibs_6_io_opinSW_0),
    .io_itrackW_0(gibs_6_io_itrackW_0),
    .io_otrackW_0(gibs_6_io_otrackW_0),
    .io_itrackN_0(gibs_6_io_itrackN_0),
    .io_otrackN_0(gibs_6_io_otrackN_0),
    .io_itrackE_0(gibs_6_io_itrackE_0),
    .io_otrackE_0(gibs_6_io_otrackE_0),
    .io_itrackS_0(gibs_6_io_itrackS_0),
    .io_otrackS_0(gibs_6_io_otrackS_0)
  );
  GIB_7 gibs_7 ( // @[CGRA.scala 333:21]
    .clock(gibs_7_clock),
    .reset(gibs_7_reset),
    .io_cfg_en(gibs_7_io_cfg_en),
    .io_cfg_addr(gibs_7_io_cfg_addr),
    .io_cfg_data(gibs_7_io_cfg_data),
    .io_ipinNW_0(gibs_7_io_ipinNW_0),
    .io_ipinNW_1(gibs_7_io_ipinNW_1),
    .io_opinNW_0(gibs_7_io_opinNW_0),
    .io_ipinNE_0(gibs_7_io_ipinNE_0),
    .io_opinNE_0(gibs_7_io_opinNE_0),
    .io_ipinSE_0(gibs_7_io_ipinSE_0),
    .io_opinSE_0(gibs_7_io_opinSE_0),
    .io_ipinSW_0(gibs_7_io_ipinSW_0),
    .io_ipinSW_1(gibs_7_io_ipinSW_1),
    .io_opinSW_0(gibs_7_io_opinSW_0),
    .io_itrackW_0(gibs_7_io_itrackW_0),
    .io_otrackW_0(gibs_7_io_otrackW_0),
    .io_itrackN_0(gibs_7_io_itrackN_0),
    .io_otrackN_0(gibs_7_io_otrackN_0),
    .io_itrackS_0(gibs_7_io_itrackS_0),
    .io_otrackS_0(gibs_7_io_otrackS_0)
  );
  GIB_8 gibs_8 ( // @[CGRA.scala 333:21]
    .clock(gibs_8_clock),
    .reset(gibs_8_reset),
    .io_cfg_en(gibs_8_io_cfg_en),
    .io_cfg_addr(gibs_8_io_cfg_addr),
    .io_cfg_data(gibs_8_io_cfg_data),
    .io_ipinNW_0(gibs_8_io_ipinNW_0),
    .io_opinNW_0(gibs_8_io_opinNW_0),
    .io_ipinNE_0(gibs_8_io_ipinNE_0),
    .io_ipinNE_1(gibs_8_io_ipinNE_1),
    .io_opinNE_0(gibs_8_io_opinNE_0),
    .io_ipinSE_0(gibs_8_io_ipinSE_0),
    .io_ipinSE_1(gibs_8_io_ipinSE_1),
    .io_opinSE_0(gibs_8_io_opinSE_0),
    .io_ipinSW_0(gibs_8_io_ipinSW_0),
    .io_opinSW_0(gibs_8_io_opinSW_0),
    .io_itrackN_0(gibs_8_io_itrackN_0),
    .io_otrackN_0(gibs_8_io_otrackN_0),
    .io_itrackE_0(gibs_8_io_itrackE_0),
    .io_otrackE_0(gibs_8_io_otrackE_0),
    .io_itrackS_0(gibs_8_io_itrackS_0),
    .io_otrackS_0(gibs_8_io_otrackS_0)
  );
  GIB_9 gibs_9 ( // @[CGRA.scala 333:21]
    .clock(gibs_9_clock),
    .reset(gibs_9_reset),
    .io_cfg_en(gibs_9_io_cfg_en),
    .io_cfg_addr(gibs_9_io_cfg_addr),
    .io_cfg_data(gibs_9_io_cfg_data),
    .io_ipinNW_0(gibs_9_io_ipinNW_0),
    .io_ipinNW_1(gibs_9_io_ipinNW_1),
    .io_opinNW_0(gibs_9_io_opinNW_0),
    .io_ipinNE_0(gibs_9_io_ipinNE_0),
    .io_ipinNE_1(gibs_9_io_ipinNE_1),
    .io_opinNE_0(gibs_9_io_opinNE_0),
    .io_ipinSE_0(gibs_9_io_ipinSE_0),
    .io_ipinSE_1(gibs_9_io_ipinSE_1),
    .io_opinSE_0(gibs_9_io_opinSE_0),
    .io_ipinSW_0(gibs_9_io_ipinSW_0),
    .io_ipinSW_1(gibs_9_io_ipinSW_1),
    .io_opinSW_0(gibs_9_io_opinSW_0),
    .io_itrackW_0(gibs_9_io_itrackW_0),
    .io_otrackW_0(gibs_9_io_otrackW_0),
    .io_itrackN_0(gibs_9_io_itrackN_0),
    .io_otrackN_0(gibs_9_io_otrackN_0),
    .io_itrackE_0(gibs_9_io_itrackE_0),
    .io_otrackE_0(gibs_9_io_otrackE_0),
    .io_itrackS_0(gibs_9_io_itrackS_0),
    .io_otrackS_0(gibs_9_io_otrackS_0)
  );
  GIB_10 gibs_10 ( // @[CGRA.scala 333:21]
    .clock(gibs_10_clock),
    .reset(gibs_10_reset),
    .io_cfg_en(gibs_10_io_cfg_en),
    .io_cfg_addr(gibs_10_io_cfg_addr),
    .io_cfg_data(gibs_10_io_cfg_data),
    .io_ipinNW_0(gibs_10_io_ipinNW_0),
    .io_ipinNW_1(gibs_10_io_ipinNW_1),
    .io_opinNW_0(gibs_10_io_opinNW_0),
    .io_ipinNE_0(gibs_10_io_ipinNE_0),
    .io_ipinNE_1(gibs_10_io_ipinNE_1),
    .io_opinNE_0(gibs_10_io_opinNE_0),
    .io_ipinSE_0(gibs_10_io_ipinSE_0),
    .io_ipinSE_1(gibs_10_io_ipinSE_1),
    .io_opinSE_0(gibs_10_io_opinSE_0),
    .io_ipinSW_0(gibs_10_io_ipinSW_0),
    .io_ipinSW_1(gibs_10_io_ipinSW_1),
    .io_opinSW_0(gibs_10_io_opinSW_0),
    .io_itrackW_0(gibs_10_io_itrackW_0),
    .io_otrackW_0(gibs_10_io_otrackW_0),
    .io_itrackN_0(gibs_10_io_itrackN_0),
    .io_otrackN_0(gibs_10_io_otrackN_0),
    .io_itrackE_0(gibs_10_io_itrackE_0),
    .io_otrackE_0(gibs_10_io_otrackE_0),
    .io_itrackS_0(gibs_10_io_itrackS_0),
    .io_otrackS_0(gibs_10_io_otrackS_0)
  );
  GIB_11 gibs_11 ( // @[CGRA.scala 333:21]
    .clock(gibs_11_clock),
    .reset(gibs_11_reset),
    .io_cfg_en(gibs_11_io_cfg_en),
    .io_cfg_addr(gibs_11_io_cfg_addr),
    .io_cfg_data(gibs_11_io_cfg_data),
    .io_ipinNW_0(gibs_11_io_ipinNW_0),
    .io_ipinNW_1(gibs_11_io_ipinNW_1),
    .io_opinNW_0(gibs_11_io_opinNW_0),
    .io_ipinNE_0(gibs_11_io_ipinNE_0),
    .io_opinNE_0(gibs_11_io_opinNE_0),
    .io_ipinSE_0(gibs_11_io_ipinSE_0),
    .io_opinSE_0(gibs_11_io_opinSE_0),
    .io_ipinSW_0(gibs_11_io_ipinSW_0),
    .io_ipinSW_1(gibs_11_io_ipinSW_1),
    .io_opinSW_0(gibs_11_io_opinSW_0),
    .io_itrackW_0(gibs_11_io_itrackW_0),
    .io_otrackW_0(gibs_11_io_otrackW_0),
    .io_itrackN_0(gibs_11_io_itrackN_0),
    .io_otrackN_0(gibs_11_io_otrackN_0),
    .io_itrackS_0(gibs_11_io_itrackS_0),
    .io_otrackS_0(gibs_11_io_otrackS_0)
  );
  GIB_12 gibs_12 ( // @[CGRA.scala 333:21]
    .clock(gibs_12_clock),
    .reset(gibs_12_reset),
    .io_cfg_en(gibs_12_io_cfg_en),
    .io_cfg_addr(gibs_12_io_cfg_addr),
    .io_cfg_data(gibs_12_io_cfg_data),
    .io_ipinNW_0(gibs_12_io_ipinNW_0),
    .io_opinNW_0(gibs_12_io_opinNW_0),
    .io_ipinNE_0(gibs_12_io_ipinNE_0),
    .io_ipinNE_1(gibs_12_io_ipinNE_1),
    .io_opinNE_0(gibs_12_io_opinNE_0),
    .io_ipinSE_0(gibs_12_io_ipinSE_0),
    .io_ipinSE_1(gibs_12_io_ipinSE_1),
    .io_opinSE_0(gibs_12_io_opinSE_0),
    .io_ipinSW_0(gibs_12_io_ipinSW_0),
    .io_opinSW_0(gibs_12_io_opinSW_0),
    .io_itrackN_0(gibs_12_io_itrackN_0),
    .io_otrackN_0(gibs_12_io_otrackN_0),
    .io_itrackE_0(gibs_12_io_itrackE_0),
    .io_otrackE_0(gibs_12_io_otrackE_0),
    .io_itrackS_0(gibs_12_io_itrackS_0),
    .io_otrackS_0(gibs_12_io_otrackS_0)
  );
  GIB_13 gibs_13 ( // @[CGRA.scala 333:21]
    .clock(gibs_13_clock),
    .reset(gibs_13_reset),
    .io_cfg_en(gibs_13_io_cfg_en),
    .io_cfg_addr(gibs_13_io_cfg_addr),
    .io_cfg_data(gibs_13_io_cfg_data),
    .io_ipinNW_0(gibs_13_io_ipinNW_0),
    .io_ipinNW_1(gibs_13_io_ipinNW_1),
    .io_opinNW_0(gibs_13_io_opinNW_0),
    .io_ipinNE_0(gibs_13_io_ipinNE_0),
    .io_ipinNE_1(gibs_13_io_ipinNE_1),
    .io_opinNE_0(gibs_13_io_opinNE_0),
    .io_ipinSE_0(gibs_13_io_ipinSE_0),
    .io_ipinSE_1(gibs_13_io_ipinSE_1),
    .io_opinSE_0(gibs_13_io_opinSE_0),
    .io_ipinSW_0(gibs_13_io_ipinSW_0),
    .io_ipinSW_1(gibs_13_io_ipinSW_1),
    .io_opinSW_0(gibs_13_io_opinSW_0),
    .io_itrackW_0(gibs_13_io_itrackW_0),
    .io_otrackW_0(gibs_13_io_otrackW_0),
    .io_itrackN_0(gibs_13_io_itrackN_0),
    .io_otrackN_0(gibs_13_io_otrackN_0),
    .io_itrackE_0(gibs_13_io_itrackE_0),
    .io_otrackE_0(gibs_13_io_otrackE_0),
    .io_itrackS_0(gibs_13_io_itrackS_0),
    .io_otrackS_0(gibs_13_io_otrackS_0)
  );
  GIB_14 gibs_14 ( // @[CGRA.scala 333:21]
    .clock(gibs_14_clock),
    .reset(gibs_14_reset),
    .io_cfg_en(gibs_14_io_cfg_en),
    .io_cfg_addr(gibs_14_io_cfg_addr),
    .io_cfg_data(gibs_14_io_cfg_data),
    .io_ipinNW_0(gibs_14_io_ipinNW_0),
    .io_ipinNW_1(gibs_14_io_ipinNW_1),
    .io_opinNW_0(gibs_14_io_opinNW_0),
    .io_ipinNE_0(gibs_14_io_ipinNE_0),
    .io_ipinNE_1(gibs_14_io_ipinNE_1),
    .io_opinNE_0(gibs_14_io_opinNE_0),
    .io_ipinSE_0(gibs_14_io_ipinSE_0),
    .io_ipinSE_1(gibs_14_io_ipinSE_1),
    .io_opinSE_0(gibs_14_io_opinSE_0),
    .io_ipinSW_0(gibs_14_io_ipinSW_0),
    .io_ipinSW_1(gibs_14_io_ipinSW_1),
    .io_opinSW_0(gibs_14_io_opinSW_0),
    .io_itrackW_0(gibs_14_io_itrackW_0),
    .io_otrackW_0(gibs_14_io_otrackW_0),
    .io_itrackN_0(gibs_14_io_itrackN_0),
    .io_otrackN_0(gibs_14_io_otrackN_0),
    .io_itrackE_0(gibs_14_io_itrackE_0),
    .io_otrackE_0(gibs_14_io_otrackE_0),
    .io_itrackS_0(gibs_14_io_itrackS_0),
    .io_otrackS_0(gibs_14_io_otrackS_0)
  );
  GIB_15 gibs_15 ( // @[CGRA.scala 333:21]
    .clock(gibs_15_clock),
    .reset(gibs_15_reset),
    .io_cfg_en(gibs_15_io_cfg_en),
    .io_cfg_addr(gibs_15_io_cfg_addr),
    .io_cfg_data(gibs_15_io_cfg_data),
    .io_ipinNW_0(gibs_15_io_ipinNW_0),
    .io_ipinNW_1(gibs_15_io_ipinNW_1),
    .io_opinNW_0(gibs_15_io_opinNW_0),
    .io_ipinNE_0(gibs_15_io_ipinNE_0),
    .io_opinNE_0(gibs_15_io_opinNE_0),
    .io_ipinSE_0(gibs_15_io_ipinSE_0),
    .io_opinSE_0(gibs_15_io_opinSE_0),
    .io_ipinSW_0(gibs_15_io_ipinSW_0),
    .io_ipinSW_1(gibs_15_io_ipinSW_1),
    .io_opinSW_0(gibs_15_io_opinSW_0),
    .io_itrackW_0(gibs_15_io_itrackW_0),
    .io_otrackW_0(gibs_15_io_otrackW_0),
    .io_itrackN_0(gibs_15_io_itrackN_0),
    .io_otrackN_0(gibs_15_io_otrackN_0),
    .io_itrackS_0(gibs_15_io_itrackS_0),
    .io_otrackS_0(gibs_15_io_otrackS_0)
  );
  GIB_16 gibs_16 ( // @[CGRA.scala 333:21]
    .clock(gibs_16_clock),
    .reset(gibs_16_reset),
    .io_cfg_en(gibs_16_io_cfg_en),
    .io_cfg_addr(gibs_16_io_cfg_addr),
    .io_cfg_data(gibs_16_io_cfg_data),
    .io_ipinNW_0(gibs_16_io_ipinNW_0),
    .io_opinNW_0(gibs_16_io_opinNW_0),
    .io_ipinNE_0(gibs_16_io_ipinNE_0),
    .io_ipinNE_1(gibs_16_io_ipinNE_1),
    .io_opinNE_0(gibs_16_io_opinNE_0),
    .io_ipinSE_0(gibs_16_io_ipinSE_0),
    .io_ipinSE_1(gibs_16_io_ipinSE_1),
    .io_opinSE_0(gibs_16_io_opinSE_0),
    .io_ipinSW_0(gibs_16_io_ipinSW_0),
    .io_opinSW_0(gibs_16_io_opinSW_0),
    .io_itrackN_0(gibs_16_io_itrackN_0),
    .io_otrackN_0(gibs_16_io_otrackN_0),
    .io_itrackE_0(gibs_16_io_itrackE_0),
    .io_otrackE_0(gibs_16_io_otrackE_0),
    .io_itrackS_0(gibs_16_io_itrackS_0),
    .io_otrackS_0(gibs_16_io_otrackS_0)
  );
  GIB_17 gibs_17 ( // @[CGRA.scala 333:21]
    .clock(gibs_17_clock),
    .reset(gibs_17_reset),
    .io_cfg_en(gibs_17_io_cfg_en),
    .io_cfg_addr(gibs_17_io_cfg_addr),
    .io_cfg_data(gibs_17_io_cfg_data),
    .io_ipinNW_0(gibs_17_io_ipinNW_0),
    .io_ipinNW_1(gibs_17_io_ipinNW_1),
    .io_opinNW_0(gibs_17_io_opinNW_0),
    .io_ipinNE_0(gibs_17_io_ipinNE_0),
    .io_ipinNE_1(gibs_17_io_ipinNE_1),
    .io_opinNE_0(gibs_17_io_opinNE_0),
    .io_ipinSE_0(gibs_17_io_ipinSE_0),
    .io_ipinSE_1(gibs_17_io_ipinSE_1),
    .io_opinSE_0(gibs_17_io_opinSE_0),
    .io_ipinSW_0(gibs_17_io_ipinSW_0),
    .io_ipinSW_1(gibs_17_io_ipinSW_1),
    .io_opinSW_0(gibs_17_io_opinSW_0),
    .io_itrackW_0(gibs_17_io_itrackW_0),
    .io_otrackW_0(gibs_17_io_otrackW_0),
    .io_itrackN_0(gibs_17_io_itrackN_0),
    .io_otrackN_0(gibs_17_io_otrackN_0),
    .io_itrackE_0(gibs_17_io_itrackE_0),
    .io_otrackE_0(gibs_17_io_otrackE_0),
    .io_itrackS_0(gibs_17_io_itrackS_0),
    .io_otrackS_0(gibs_17_io_otrackS_0)
  );
  GIB_18 gibs_18 ( // @[CGRA.scala 333:21]
    .clock(gibs_18_clock),
    .reset(gibs_18_reset),
    .io_cfg_en(gibs_18_io_cfg_en),
    .io_cfg_addr(gibs_18_io_cfg_addr),
    .io_cfg_data(gibs_18_io_cfg_data),
    .io_ipinNW_0(gibs_18_io_ipinNW_0),
    .io_ipinNW_1(gibs_18_io_ipinNW_1),
    .io_opinNW_0(gibs_18_io_opinNW_0),
    .io_ipinNE_0(gibs_18_io_ipinNE_0),
    .io_ipinNE_1(gibs_18_io_ipinNE_1),
    .io_opinNE_0(gibs_18_io_opinNE_0),
    .io_ipinSE_0(gibs_18_io_ipinSE_0),
    .io_ipinSE_1(gibs_18_io_ipinSE_1),
    .io_opinSE_0(gibs_18_io_opinSE_0),
    .io_ipinSW_0(gibs_18_io_ipinSW_0),
    .io_ipinSW_1(gibs_18_io_ipinSW_1),
    .io_opinSW_0(gibs_18_io_opinSW_0),
    .io_itrackW_0(gibs_18_io_itrackW_0),
    .io_otrackW_0(gibs_18_io_otrackW_0),
    .io_itrackN_0(gibs_18_io_itrackN_0),
    .io_otrackN_0(gibs_18_io_otrackN_0),
    .io_itrackE_0(gibs_18_io_itrackE_0),
    .io_otrackE_0(gibs_18_io_otrackE_0),
    .io_itrackS_0(gibs_18_io_itrackS_0),
    .io_otrackS_0(gibs_18_io_otrackS_0)
  );
  GIB_19 gibs_19 ( // @[CGRA.scala 333:21]
    .clock(gibs_19_clock),
    .reset(gibs_19_reset),
    .io_cfg_en(gibs_19_io_cfg_en),
    .io_cfg_addr(gibs_19_io_cfg_addr),
    .io_cfg_data(gibs_19_io_cfg_data),
    .io_ipinNW_0(gibs_19_io_ipinNW_0),
    .io_ipinNW_1(gibs_19_io_ipinNW_1),
    .io_opinNW_0(gibs_19_io_opinNW_0),
    .io_ipinNE_0(gibs_19_io_ipinNE_0),
    .io_opinNE_0(gibs_19_io_opinNE_0),
    .io_ipinSE_0(gibs_19_io_ipinSE_0),
    .io_opinSE_0(gibs_19_io_opinSE_0),
    .io_ipinSW_0(gibs_19_io_ipinSW_0),
    .io_ipinSW_1(gibs_19_io_ipinSW_1),
    .io_opinSW_0(gibs_19_io_opinSW_0),
    .io_itrackW_0(gibs_19_io_itrackW_0),
    .io_otrackW_0(gibs_19_io_otrackW_0),
    .io_itrackN_0(gibs_19_io_itrackN_0),
    .io_otrackN_0(gibs_19_io_otrackN_0),
    .io_itrackS_0(gibs_19_io_itrackS_0),
    .io_otrackS_0(gibs_19_io_otrackS_0)
  );
  GIB_20 gibs_20 ( // @[CGRA.scala 333:21]
    .clock(gibs_20_clock),
    .reset(gibs_20_reset),
    .io_cfg_en(gibs_20_io_cfg_en),
    .io_cfg_addr(gibs_20_io_cfg_addr),
    .io_cfg_data(gibs_20_io_cfg_data),
    .io_ipinNW_0(gibs_20_io_ipinNW_0),
    .io_opinNW_0(gibs_20_io_opinNW_0),
    .io_ipinNE_0(gibs_20_io_ipinNE_0),
    .io_ipinNE_1(gibs_20_io_ipinNE_1),
    .io_opinNE_0(gibs_20_io_opinNE_0),
    .io_ipinSE_0(gibs_20_io_ipinSE_0),
    .io_ipinSE_1(gibs_20_io_ipinSE_1),
    .io_opinSE_0(gibs_20_io_opinSE_0),
    .io_ipinSW_0(gibs_20_io_ipinSW_0),
    .io_opinSW_0(gibs_20_io_opinSW_0),
    .io_itrackN_0(gibs_20_io_itrackN_0),
    .io_otrackN_0(gibs_20_io_otrackN_0),
    .io_itrackE_0(gibs_20_io_itrackE_0),
    .io_otrackE_0(gibs_20_io_otrackE_0),
    .io_itrackS_0(gibs_20_io_itrackS_0),
    .io_otrackS_0(gibs_20_io_otrackS_0)
  );
  GIB_21 gibs_21 ( // @[CGRA.scala 333:21]
    .clock(gibs_21_clock),
    .reset(gibs_21_reset),
    .io_cfg_en(gibs_21_io_cfg_en),
    .io_cfg_addr(gibs_21_io_cfg_addr),
    .io_cfg_data(gibs_21_io_cfg_data),
    .io_ipinNW_0(gibs_21_io_ipinNW_0),
    .io_ipinNW_1(gibs_21_io_ipinNW_1),
    .io_opinNW_0(gibs_21_io_opinNW_0),
    .io_ipinNE_0(gibs_21_io_ipinNE_0),
    .io_ipinNE_1(gibs_21_io_ipinNE_1),
    .io_opinNE_0(gibs_21_io_opinNE_0),
    .io_ipinSE_0(gibs_21_io_ipinSE_0),
    .io_ipinSE_1(gibs_21_io_ipinSE_1),
    .io_opinSE_0(gibs_21_io_opinSE_0),
    .io_ipinSW_0(gibs_21_io_ipinSW_0),
    .io_ipinSW_1(gibs_21_io_ipinSW_1),
    .io_opinSW_0(gibs_21_io_opinSW_0),
    .io_itrackW_0(gibs_21_io_itrackW_0),
    .io_otrackW_0(gibs_21_io_otrackW_0),
    .io_itrackN_0(gibs_21_io_itrackN_0),
    .io_otrackN_0(gibs_21_io_otrackN_0),
    .io_itrackE_0(gibs_21_io_itrackE_0),
    .io_otrackE_0(gibs_21_io_otrackE_0),
    .io_itrackS_0(gibs_21_io_itrackS_0),
    .io_otrackS_0(gibs_21_io_otrackS_0)
  );
  GIB_22 gibs_22 ( // @[CGRA.scala 333:21]
    .clock(gibs_22_clock),
    .reset(gibs_22_reset),
    .io_cfg_en(gibs_22_io_cfg_en),
    .io_cfg_addr(gibs_22_io_cfg_addr),
    .io_cfg_data(gibs_22_io_cfg_data),
    .io_ipinNW_0(gibs_22_io_ipinNW_0),
    .io_ipinNW_1(gibs_22_io_ipinNW_1),
    .io_opinNW_0(gibs_22_io_opinNW_0),
    .io_ipinNE_0(gibs_22_io_ipinNE_0),
    .io_ipinNE_1(gibs_22_io_ipinNE_1),
    .io_opinNE_0(gibs_22_io_opinNE_0),
    .io_ipinSE_0(gibs_22_io_ipinSE_0),
    .io_ipinSE_1(gibs_22_io_ipinSE_1),
    .io_opinSE_0(gibs_22_io_opinSE_0),
    .io_ipinSW_0(gibs_22_io_ipinSW_0),
    .io_ipinSW_1(gibs_22_io_ipinSW_1),
    .io_opinSW_0(gibs_22_io_opinSW_0),
    .io_itrackW_0(gibs_22_io_itrackW_0),
    .io_otrackW_0(gibs_22_io_otrackW_0),
    .io_itrackN_0(gibs_22_io_itrackN_0),
    .io_otrackN_0(gibs_22_io_otrackN_0),
    .io_itrackE_0(gibs_22_io_itrackE_0),
    .io_otrackE_0(gibs_22_io_otrackE_0),
    .io_itrackS_0(gibs_22_io_itrackS_0),
    .io_otrackS_0(gibs_22_io_otrackS_0)
  );
  GIB_23 gibs_23 ( // @[CGRA.scala 333:21]
    .clock(gibs_23_clock),
    .reset(gibs_23_reset),
    .io_cfg_en(gibs_23_io_cfg_en),
    .io_cfg_addr(gibs_23_io_cfg_addr),
    .io_cfg_data(gibs_23_io_cfg_data),
    .io_ipinNW_0(gibs_23_io_ipinNW_0),
    .io_ipinNW_1(gibs_23_io_ipinNW_1),
    .io_opinNW_0(gibs_23_io_opinNW_0),
    .io_ipinNE_0(gibs_23_io_ipinNE_0),
    .io_opinNE_0(gibs_23_io_opinNE_0),
    .io_ipinSE_0(gibs_23_io_ipinSE_0),
    .io_opinSE_0(gibs_23_io_opinSE_0),
    .io_ipinSW_0(gibs_23_io_ipinSW_0),
    .io_ipinSW_1(gibs_23_io_ipinSW_1),
    .io_opinSW_0(gibs_23_io_opinSW_0),
    .io_itrackW_0(gibs_23_io_itrackW_0),
    .io_otrackW_0(gibs_23_io_otrackW_0),
    .io_itrackN_0(gibs_23_io_itrackN_0),
    .io_otrackN_0(gibs_23_io_otrackN_0),
    .io_itrackS_0(gibs_23_io_itrackS_0),
    .io_otrackS_0(gibs_23_io_otrackS_0)
  );
  GIB_24 gibs_24 ( // @[CGRA.scala 333:21]
    .clock(gibs_24_clock),
    .reset(gibs_24_reset),
    .io_cfg_en(gibs_24_io_cfg_en),
    .io_cfg_addr(gibs_24_io_cfg_addr),
    .io_cfg_data(gibs_24_io_cfg_data),
    .io_ipinNW_0(gibs_24_io_ipinNW_0),
    .io_opinNW_0(gibs_24_io_opinNW_0),
    .io_ipinNE_0(gibs_24_io_ipinNE_0),
    .io_ipinNE_1(gibs_24_io_ipinNE_1),
    .io_opinNE_0(gibs_24_io_opinNE_0),
    .io_ipinSE_0(gibs_24_io_ipinSE_0),
    .io_ipinSE_1(gibs_24_io_ipinSE_1),
    .io_opinSE_0(gibs_24_io_opinSE_0),
    .io_ipinSW_0(gibs_24_io_ipinSW_0),
    .io_opinSW_0(gibs_24_io_opinSW_0),
    .io_itrackN_0(gibs_24_io_itrackN_0),
    .io_otrackN_0(gibs_24_io_otrackN_0),
    .io_itrackE_0(gibs_24_io_itrackE_0),
    .io_otrackE_0(gibs_24_io_otrackE_0),
    .io_itrackS_0(gibs_24_io_itrackS_0),
    .io_otrackS_0(gibs_24_io_otrackS_0)
  );
  GIB_25 gibs_25 ( // @[CGRA.scala 333:21]
    .clock(gibs_25_clock),
    .reset(gibs_25_reset),
    .io_cfg_en(gibs_25_io_cfg_en),
    .io_cfg_addr(gibs_25_io_cfg_addr),
    .io_cfg_data(gibs_25_io_cfg_data),
    .io_ipinNW_0(gibs_25_io_ipinNW_0),
    .io_ipinNW_1(gibs_25_io_ipinNW_1),
    .io_opinNW_0(gibs_25_io_opinNW_0),
    .io_ipinNE_0(gibs_25_io_ipinNE_0),
    .io_ipinNE_1(gibs_25_io_ipinNE_1),
    .io_opinNE_0(gibs_25_io_opinNE_0),
    .io_ipinSE_0(gibs_25_io_ipinSE_0),
    .io_ipinSE_1(gibs_25_io_ipinSE_1),
    .io_opinSE_0(gibs_25_io_opinSE_0),
    .io_ipinSW_0(gibs_25_io_ipinSW_0),
    .io_ipinSW_1(gibs_25_io_ipinSW_1),
    .io_opinSW_0(gibs_25_io_opinSW_0),
    .io_itrackW_0(gibs_25_io_itrackW_0),
    .io_otrackW_0(gibs_25_io_otrackW_0),
    .io_itrackN_0(gibs_25_io_itrackN_0),
    .io_otrackN_0(gibs_25_io_otrackN_0),
    .io_itrackE_0(gibs_25_io_itrackE_0),
    .io_otrackE_0(gibs_25_io_otrackE_0),
    .io_itrackS_0(gibs_25_io_itrackS_0),
    .io_otrackS_0(gibs_25_io_otrackS_0)
  );
  GIB_26 gibs_26 ( // @[CGRA.scala 333:21]
    .clock(gibs_26_clock),
    .reset(gibs_26_reset),
    .io_cfg_en(gibs_26_io_cfg_en),
    .io_cfg_addr(gibs_26_io_cfg_addr),
    .io_cfg_data(gibs_26_io_cfg_data),
    .io_ipinNW_0(gibs_26_io_ipinNW_0),
    .io_ipinNW_1(gibs_26_io_ipinNW_1),
    .io_opinNW_0(gibs_26_io_opinNW_0),
    .io_ipinNE_0(gibs_26_io_ipinNE_0),
    .io_ipinNE_1(gibs_26_io_ipinNE_1),
    .io_opinNE_0(gibs_26_io_opinNE_0),
    .io_ipinSE_0(gibs_26_io_ipinSE_0),
    .io_ipinSE_1(gibs_26_io_ipinSE_1),
    .io_opinSE_0(gibs_26_io_opinSE_0),
    .io_ipinSW_0(gibs_26_io_ipinSW_0),
    .io_ipinSW_1(gibs_26_io_ipinSW_1),
    .io_opinSW_0(gibs_26_io_opinSW_0),
    .io_itrackW_0(gibs_26_io_itrackW_0),
    .io_otrackW_0(gibs_26_io_otrackW_0),
    .io_itrackN_0(gibs_26_io_itrackN_0),
    .io_otrackN_0(gibs_26_io_otrackN_0),
    .io_itrackE_0(gibs_26_io_itrackE_0),
    .io_otrackE_0(gibs_26_io_otrackE_0),
    .io_itrackS_0(gibs_26_io_itrackS_0),
    .io_otrackS_0(gibs_26_io_otrackS_0)
  );
  GIB_27 gibs_27 ( // @[CGRA.scala 333:21]
    .clock(gibs_27_clock),
    .reset(gibs_27_reset),
    .io_cfg_en(gibs_27_io_cfg_en),
    .io_cfg_addr(gibs_27_io_cfg_addr),
    .io_cfg_data(gibs_27_io_cfg_data),
    .io_ipinNW_0(gibs_27_io_ipinNW_0),
    .io_ipinNW_1(gibs_27_io_ipinNW_1),
    .io_opinNW_0(gibs_27_io_opinNW_0),
    .io_ipinNE_0(gibs_27_io_ipinNE_0),
    .io_opinNE_0(gibs_27_io_opinNE_0),
    .io_ipinSE_0(gibs_27_io_ipinSE_0),
    .io_opinSE_0(gibs_27_io_opinSE_0),
    .io_ipinSW_0(gibs_27_io_ipinSW_0),
    .io_ipinSW_1(gibs_27_io_ipinSW_1),
    .io_opinSW_0(gibs_27_io_opinSW_0),
    .io_itrackW_0(gibs_27_io_itrackW_0),
    .io_otrackW_0(gibs_27_io_otrackW_0),
    .io_itrackN_0(gibs_27_io_itrackN_0),
    .io_otrackN_0(gibs_27_io_otrackN_0),
    .io_itrackS_0(gibs_27_io_itrackS_0),
    .io_otrackS_0(gibs_27_io_otrackS_0)
  );
  GIB_28 gibs_28 ( // @[CGRA.scala 333:21]
    .clock(gibs_28_clock),
    .reset(gibs_28_reset),
    .io_cfg_en(gibs_28_io_cfg_en),
    .io_cfg_addr(gibs_28_io_cfg_addr),
    .io_cfg_data(gibs_28_io_cfg_data),
    .io_ipinNW_0(gibs_28_io_ipinNW_0),
    .io_opinNW_0(gibs_28_io_opinNW_0),
    .io_ipinNE_0(gibs_28_io_ipinNE_0),
    .io_ipinNE_1(gibs_28_io_ipinNE_1),
    .io_opinNE_0(gibs_28_io_opinNE_0),
    .io_ipinSE_0(gibs_28_io_ipinSE_0),
    .io_ipinSE_1(gibs_28_io_ipinSE_1),
    .io_opinSE_0(gibs_28_io_opinSE_0),
    .io_ipinSW_0(gibs_28_io_ipinSW_0),
    .io_opinSW_0(gibs_28_io_opinSW_0),
    .io_itrackN_0(gibs_28_io_itrackN_0),
    .io_otrackN_0(gibs_28_io_otrackN_0),
    .io_itrackE_0(gibs_28_io_itrackE_0),
    .io_otrackE_0(gibs_28_io_otrackE_0),
    .io_itrackS_0(gibs_28_io_itrackS_0),
    .io_otrackS_0(gibs_28_io_otrackS_0)
  );
  GIB_29 gibs_29 ( // @[CGRA.scala 333:21]
    .clock(gibs_29_clock),
    .reset(gibs_29_reset),
    .io_cfg_en(gibs_29_io_cfg_en),
    .io_cfg_addr(gibs_29_io_cfg_addr),
    .io_cfg_data(gibs_29_io_cfg_data),
    .io_ipinNW_0(gibs_29_io_ipinNW_0),
    .io_ipinNW_1(gibs_29_io_ipinNW_1),
    .io_opinNW_0(gibs_29_io_opinNW_0),
    .io_ipinNE_0(gibs_29_io_ipinNE_0),
    .io_ipinNE_1(gibs_29_io_ipinNE_1),
    .io_opinNE_0(gibs_29_io_opinNE_0),
    .io_ipinSE_0(gibs_29_io_ipinSE_0),
    .io_ipinSE_1(gibs_29_io_ipinSE_1),
    .io_opinSE_0(gibs_29_io_opinSE_0),
    .io_ipinSW_0(gibs_29_io_ipinSW_0),
    .io_ipinSW_1(gibs_29_io_ipinSW_1),
    .io_opinSW_0(gibs_29_io_opinSW_0),
    .io_itrackW_0(gibs_29_io_itrackW_0),
    .io_otrackW_0(gibs_29_io_otrackW_0),
    .io_itrackN_0(gibs_29_io_itrackN_0),
    .io_otrackN_0(gibs_29_io_otrackN_0),
    .io_itrackE_0(gibs_29_io_itrackE_0),
    .io_otrackE_0(gibs_29_io_otrackE_0),
    .io_itrackS_0(gibs_29_io_itrackS_0),
    .io_otrackS_0(gibs_29_io_otrackS_0)
  );
  GIB_30 gibs_30 ( // @[CGRA.scala 333:21]
    .clock(gibs_30_clock),
    .reset(gibs_30_reset),
    .io_cfg_en(gibs_30_io_cfg_en),
    .io_cfg_addr(gibs_30_io_cfg_addr),
    .io_cfg_data(gibs_30_io_cfg_data),
    .io_ipinNW_0(gibs_30_io_ipinNW_0),
    .io_ipinNW_1(gibs_30_io_ipinNW_1),
    .io_opinNW_0(gibs_30_io_opinNW_0),
    .io_ipinNE_0(gibs_30_io_ipinNE_0),
    .io_ipinNE_1(gibs_30_io_ipinNE_1),
    .io_opinNE_0(gibs_30_io_opinNE_0),
    .io_ipinSE_0(gibs_30_io_ipinSE_0),
    .io_ipinSE_1(gibs_30_io_ipinSE_1),
    .io_opinSE_0(gibs_30_io_opinSE_0),
    .io_ipinSW_0(gibs_30_io_ipinSW_0),
    .io_ipinSW_1(gibs_30_io_ipinSW_1),
    .io_opinSW_0(gibs_30_io_opinSW_0),
    .io_itrackW_0(gibs_30_io_itrackW_0),
    .io_otrackW_0(gibs_30_io_otrackW_0),
    .io_itrackN_0(gibs_30_io_itrackN_0),
    .io_otrackN_0(gibs_30_io_otrackN_0),
    .io_itrackE_0(gibs_30_io_itrackE_0),
    .io_otrackE_0(gibs_30_io_otrackE_0),
    .io_itrackS_0(gibs_30_io_itrackS_0),
    .io_otrackS_0(gibs_30_io_otrackS_0)
  );
  GIB_31 gibs_31 ( // @[CGRA.scala 333:21]
    .clock(gibs_31_clock),
    .reset(gibs_31_reset),
    .io_cfg_en(gibs_31_io_cfg_en),
    .io_cfg_addr(gibs_31_io_cfg_addr),
    .io_cfg_data(gibs_31_io_cfg_data),
    .io_ipinNW_0(gibs_31_io_ipinNW_0),
    .io_ipinNW_1(gibs_31_io_ipinNW_1),
    .io_opinNW_0(gibs_31_io_opinNW_0),
    .io_ipinNE_0(gibs_31_io_ipinNE_0),
    .io_opinNE_0(gibs_31_io_opinNE_0),
    .io_ipinSE_0(gibs_31_io_ipinSE_0),
    .io_opinSE_0(gibs_31_io_opinSE_0),
    .io_ipinSW_0(gibs_31_io_ipinSW_0),
    .io_ipinSW_1(gibs_31_io_ipinSW_1),
    .io_opinSW_0(gibs_31_io_opinSW_0),
    .io_itrackW_0(gibs_31_io_itrackW_0),
    .io_otrackW_0(gibs_31_io_otrackW_0),
    .io_itrackN_0(gibs_31_io_itrackN_0),
    .io_otrackN_0(gibs_31_io_otrackN_0),
    .io_itrackS_0(gibs_31_io_itrackS_0),
    .io_otrackS_0(gibs_31_io_otrackS_0)
  );
  GIB_32 gibs_32 ( // @[CGRA.scala 333:21]
    .clock(gibs_32_clock),
    .reset(gibs_32_reset),
    .io_cfg_en(gibs_32_io_cfg_en),
    .io_cfg_addr(gibs_32_io_cfg_addr),
    .io_cfg_data(gibs_32_io_cfg_data),
    .io_ipinNW_0(gibs_32_io_ipinNW_0),
    .io_opinNW_0(gibs_32_io_opinNW_0),
    .io_ipinNE_0(gibs_32_io_ipinNE_0),
    .io_ipinNE_1(gibs_32_io_ipinNE_1),
    .io_opinNE_0(gibs_32_io_opinNE_0),
    .io_ipinSE_0(gibs_32_io_ipinSE_0),
    .io_ipinSE_1(gibs_32_io_ipinSE_1),
    .io_opinSE_0(gibs_32_io_opinSE_0),
    .io_ipinSW_0(gibs_32_io_ipinSW_0),
    .io_opinSW_0(gibs_32_io_opinSW_0),
    .io_itrackN_0(gibs_32_io_itrackN_0),
    .io_otrackN_0(gibs_32_io_otrackN_0),
    .io_itrackE_0(gibs_32_io_itrackE_0),
    .io_otrackE_0(gibs_32_io_otrackE_0),
    .io_itrackS_0(gibs_32_io_itrackS_0),
    .io_otrackS_0(gibs_32_io_otrackS_0)
  );
  GIB_33 gibs_33 ( // @[CGRA.scala 333:21]
    .clock(gibs_33_clock),
    .reset(gibs_33_reset),
    .io_cfg_en(gibs_33_io_cfg_en),
    .io_cfg_addr(gibs_33_io_cfg_addr),
    .io_cfg_data(gibs_33_io_cfg_data),
    .io_ipinNW_0(gibs_33_io_ipinNW_0),
    .io_ipinNW_1(gibs_33_io_ipinNW_1),
    .io_opinNW_0(gibs_33_io_opinNW_0),
    .io_ipinNE_0(gibs_33_io_ipinNE_0),
    .io_ipinNE_1(gibs_33_io_ipinNE_1),
    .io_opinNE_0(gibs_33_io_opinNE_0),
    .io_ipinSE_0(gibs_33_io_ipinSE_0),
    .io_ipinSE_1(gibs_33_io_ipinSE_1),
    .io_opinSE_0(gibs_33_io_opinSE_0),
    .io_ipinSW_0(gibs_33_io_ipinSW_0),
    .io_ipinSW_1(gibs_33_io_ipinSW_1),
    .io_opinSW_0(gibs_33_io_opinSW_0),
    .io_itrackW_0(gibs_33_io_itrackW_0),
    .io_otrackW_0(gibs_33_io_otrackW_0),
    .io_itrackN_0(gibs_33_io_itrackN_0),
    .io_otrackN_0(gibs_33_io_otrackN_0),
    .io_itrackE_0(gibs_33_io_itrackE_0),
    .io_otrackE_0(gibs_33_io_otrackE_0),
    .io_itrackS_0(gibs_33_io_itrackS_0),
    .io_otrackS_0(gibs_33_io_otrackS_0)
  );
  GIB_34 gibs_34 ( // @[CGRA.scala 333:21]
    .clock(gibs_34_clock),
    .reset(gibs_34_reset),
    .io_cfg_en(gibs_34_io_cfg_en),
    .io_cfg_addr(gibs_34_io_cfg_addr),
    .io_cfg_data(gibs_34_io_cfg_data),
    .io_ipinNW_0(gibs_34_io_ipinNW_0),
    .io_ipinNW_1(gibs_34_io_ipinNW_1),
    .io_opinNW_0(gibs_34_io_opinNW_0),
    .io_ipinNE_0(gibs_34_io_ipinNE_0),
    .io_ipinNE_1(gibs_34_io_ipinNE_1),
    .io_opinNE_0(gibs_34_io_opinNE_0),
    .io_ipinSE_0(gibs_34_io_ipinSE_0),
    .io_ipinSE_1(gibs_34_io_ipinSE_1),
    .io_opinSE_0(gibs_34_io_opinSE_0),
    .io_ipinSW_0(gibs_34_io_ipinSW_0),
    .io_ipinSW_1(gibs_34_io_ipinSW_1),
    .io_opinSW_0(gibs_34_io_opinSW_0),
    .io_itrackW_0(gibs_34_io_itrackW_0),
    .io_otrackW_0(gibs_34_io_otrackW_0),
    .io_itrackN_0(gibs_34_io_itrackN_0),
    .io_otrackN_0(gibs_34_io_otrackN_0),
    .io_itrackE_0(gibs_34_io_itrackE_0),
    .io_otrackE_0(gibs_34_io_otrackE_0),
    .io_itrackS_0(gibs_34_io_itrackS_0),
    .io_otrackS_0(gibs_34_io_otrackS_0)
  );
  GIB_35 gibs_35 ( // @[CGRA.scala 333:21]
    .clock(gibs_35_clock),
    .reset(gibs_35_reset),
    .io_cfg_en(gibs_35_io_cfg_en),
    .io_cfg_addr(gibs_35_io_cfg_addr),
    .io_cfg_data(gibs_35_io_cfg_data),
    .io_ipinNW_0(gibs_35_io_ipinNW_0),
    .io_ipinNW_1(gibs_35_io_ipinNW_1),
    .io_opinNW_0(gibs_35_io_opinNW_0),
    .io_ipinNE_0(gibs_35_io_ipinNE_0),
    .io_opinNE_0(gibs_35_io_opinNE_0),
    .io_ipinSE_0(gibs_35_io_ipinSE_0),
    .io_opinSE_0(gibs_35_io_opinSE_0),
    .io_ipinSW_0(gibs_35_io_ipinSW_0),
    .io_ipinSW_1(gibs_35_io_ipinSW_1),
    .io_opinSW_0(gibs_35_io_opinSW_0),
    .io_itrackW_0(gibs_35_io_itrackW_0),
    .io_otrackW_0(gibs_35_io_otrackW_0),
    .io_itrackN_0(gibs_35_io_itrackN_0),
    .io_otrackN_0(gibs_35_io_otrackN_0),
    .io_itrackS_0(gibs_35_io_itrackS_0),
    .io_otrackS_0(gibs_35_io_otrackS_0)
  );
  GIB_36 gibs_36 ( // @[CGRA.scala 333:21]
    .clock(gibs_36_clock),
    .reset(gibs_36_reset),
    .io_cfg_en(gibs_36_io_cfg_en),
    .io_cfg_addr(gibs_36_io_cfg_addr),
    .io_cfg_data(gibs_36_io_cfg_data),
    .io_ipinNW_0(gibs_36_io_ipinNW_0),
    .io_opinNW_0(gibs_36_io_opinNW_0),
    .io_ipinNE_0(gibs_36_io_ipinNE_0),
    .io_ipinNE_1(gibs_36_io_ipinNE_1),
    .io_opinNE_0(gibs_36_io_opinNE_0),
    .io_ipinSE_0(gibs_36_io_ipinSE_0),
    .io_ipinSE_1(gibs_36_io_ipinSE_1),
    .io_opinSE_0(gibs_36_io_opinSE_0),
    .io_ipinSW_0(gibs_36_io_ipinSW_0),
    .io_opinSW_0(gibs_36_io_opinSW_0),
    .io_itrackN_0(gibs_36_io_itrackN_0),
    .io_otrackN_0(gibs_36_io_otrackN_0),
    .io_itrackE_0(gibs_36_io_itrackE_0),
    .io_otrackE_0(gibs_36_io_otrackE_0),
    .io_itrackS_0(gibs_36_io_itrackS_0),
    .io_otrackS_0(gibs_36_io_otrackS_0)
  );
  GIB_37 gibs_37 ( // @[CGRA.scala 333:21]
    .clock(gibs_37_clock),
    .reset(gibs_37_reset),
    .io_cfg_en(gibs_37_io_cfg_en),
    .io_cfg_addr(gibs_37_io_cfg_addr),
    .io_cfg_data(gibs_37_io_cfg_data),
    .io_ipinNW_0(gibs_37_io_ipinNW_0),
    .io_ipinNW_1(gibs_37_io_ipinNW_1),
    .io_opinNW_0(gibs_37_io_opinNW_0),
    .io_ipinNE_0(gibs_37_io_ipinNE_0),
    .io_ipinNE_1(gibs_37_io_ipinNE_1),
    .io_opinNE_0(gibs_37_io_opinNE_0),
    .io_ipinSE_0(gibs_37_io_ipinSE_0),
    .io_ipinSE_1(gibs_37_io_ipinSE_1),
    .io_opinSE_0(gibs_37_io_opinSE_0),
    .io_ipinSW_0(gibs_37_io_ipinSW_0),
    .io_ipinSW_1(gibs_37_io_ipinSW_1),
    .io_opinSW_0(gibs_37_io_opinSW_0),
    .io_itrackW_0(gibs_37_io_itrackW_0),
    .io_otrackW_0(gibs_37_io_otrackW_0),
    .io_itrackN_0(gibs_37_io_itrackN_0),
    .io_otrackN_0(gibs_37_io_otrackN_0),
    .io_itrackE_0(gibs_37_io_itrackE_0),
    .io_otrackE_0(gibs_37_io_otrackE_0),
    .io_itrackS_0(gibs_37_io_itrackS_0),
    .io_otrackS_0(gibs_37_io_otrackS_0)
  );
  GIB_38 gibs_38 ( // @[CGRA.scala 333:21]
    .clock(gibs_38_clock),
    .reset(gibs_38_reset),
    .io_cfg_en(gibs_38_io_cfg_en),
    .io_cfg_addr(gibs_38_io_cfg_addr),
    .io_cfg_data(gibs_38_io_cfg_data),
    .io_ipinNW_0(gibs_38_io_ipinNW_0),
    .io_ipinNW_1(gibs_38_io_ipinNW_1),
    .io_opinNW_0(gibs_38_io_opinNW_0),
    .io_ipinNE_0(gibs_38_io_ipinNE_0),
    .io_ipinNE_1(gibs_38_io_ipinNE_1),
    .io_opinNE_0(gibs_38_io_opinNE_0),
    .io_ipinSE_0(gibs_38_io_ipinSE_0),
    .io_ipinSE_1(gibs_38_io_ipinSE_1),
    .io_opinSE_0(gibs_38_io_opinSE_0),
    .io_ipinSW_0(gibs_38_io_ipinSW_0),
    .io_ipinSW_1(gibs_38_io_ipinSW_1),
    .io_opinSW_0(gibs_38_io_opinSW_0),
    .io_itrackW_0(gibs_38_io_itrackW_0),
    .io_otrackW_0(gibs_38_io_otrackW_0),
    .io_itrackN_0(gibs_38_io_itrackN_0),
    .io_otrackN_0(gibs_38_io_otrackN_0),
    .io_itrackE_0(gibs_38_io_itrackE_0),
    .io_otrackE_0(gibs_38_io_otrackE_0),
    .io_itrackS_0(gibs_38_io_itrackS_0),
    .io_otrackS_0(gibs_38_io_otrackS_0)
  );
  GIB_39 gibs_39 ( // @[CGRA.scala 333:21]
    .clock(gibs_39_clock),
    .reset(gibs_39_reset),
    .io_cfg_en(gibs_39_io_cfg_en),
    .io_cfg_addr(gibs_39_io_cfg_addr),
    .io_cfg_data(gibs_39_io_cfg_data),
    .io_ipinNW_0(gibs_39_io_ipinNW_0),
    .io_ipinNW_1(gibs_39_io_ipinNW_1),
    .io_opinNW_0(gibs_39_io_opinNW_0),
    .io_ipinNE_0(gibs_39_io_ipinNE_0),
    .io_opinNE_0(gibs_39_io_opinNE_0),
    .io_ipinSE_0(gibs_39_io_ipinSE_0),
    .io_opinSE_0(gibs_39_io_opinSE_0),
    .io_ipinSW_0(gibs_39_io_ipinSW_0),
    .io_ipinSW_1(gibs_39_io_ipinSW_1),
    .io_opinSW_0(gibs_39_io_opinSW_0),
    .io_itrackW_0(gibs_39_io_itrackW_0),
    .io_otrackW_0(gibs_39_io_otrackW_0),
    .io_itrackN_0(gibs_39_io_itrackN_0),
    .io_otrackN_0(gibs_39_io_otrackN_0),
    .io_itrackS_0(gibs_39_io_itrackS_0),
    .io_otrackS_0(gibs_39_io_otrackS_0)
  );
  GIB_40 gibs_40 ( // @[CGRA.scala 333:21]
    .clock(gibs_40_clock),
    .reset(gibs_40_reset),
    .io_cfg_en(gibs_40_io_cfg_en),
    .io_cfg_addr(gibs_40_io_cfg_addr),
    .io_cfg_data(gibs_40_io_cfg_data),
    .io_ipinNW_0(gibs_40_io_ipinNW_0),
    .io_opinNW_0(gibs_40_io_opinNW_0),
    .io_ipinNE_0(gibs_40_io_ipinNE_0),
    .io_ipinNE_1(gibs_40_io_ipinNE_1),
    .io_opinNE_0(gibs_40_io_opinNE_0),
    .io_ipinSE_0(gibs_40_io_ipinSE_0),
    .io_ipinSE_1(gibs_40_io_ipinSE_1),
    .io_opinSE_0(gibs_40_io_opinSE_0),
    .io_ipinSW_0(gibs_40_io_ipinSW_0),
    .io_opinSW_0(gibs_40_io_opinSW_0),
    .io_itrackN_0(gibs_40_io_itrackN_0),
    .io_otrackN_0(gibs_40_io_otrackN_0),
    .io_itrackE_0(gibs_40_io_itrackE_0),
    .io_otrackE_0(gibs_40_io_otrackE_0),
    .io_itrackS_0(gibs_40_io_itrackS_0),
    .io_otrackS_0(gibs_40_io_otrackS_0)
  );
  GIB_41 gibs_41 ( // @[CGRA.scala 333:21]
    .clock(gibs_41_clock),
    .reset(gibs_41_reset),
    .io_cfg_en(gibs_41_io_cfg_en),
    .io_cfg_addr(gibs_41_io_cfg_addr),
    .io_cfg_data(gibs_41_io_cfg_data),
    .io_ipinNW_0(gibs_41_io_ipinNW_0),
    .io_ipinNW_1(gibs_41_io_ipinNW_1),
    .io_opinNW_0(gibs_41_io_opinNW_0),
    .io_ipinNE_0(gibs_41_io_ipinNE_0),
    .io_ipinNE_1(gibs_41_io_ipinNE_1),
    .io_opinNE_0(gibs_41_io_opinNE_0),
    .io_ipinSE_0(gibs_41_io_ipinSE_0),
    .io_ipinSE_1(gibs_41_io_ipinSE_1),
    .io_opinSE_0(gibs_41_io_opinSE_0),
    .io_ipinSW_0(gibs_41_io_ipinSW_0),
    .io_ipinSW_1(gibs_41_io_ipinSW_1),
    .io_opinSW_0(gibs_41_io_opinSW_0),
    .io_itrackW_0(gibs_41_io_itrackW_0),
    .io_otrackW_0(gibs_41_io_otrackW_0),
    .io_itrackN_0(gibs_41_io_itrackN_0),
    .io_otrackN_0(gibs_41_io_otrackN_0),
    .io_itrackE_0(gibs_41_io_itrackE_0),
    .io_otrackE_0(gibs_41_io_otrackE_0),
    .io_itrackS_0(gibs_41_io_itrackS_0),
    .io_otrackS_0(gibs_41_io_otrackS_0)
  );
  GIB_42 gibs_42 ( // @[CGRA.scala 333:21]
    .clock(gibs_42_clock),
    .reset(gibs_42_reset),
    .io_cfg_en(gibs_42_io_cfg_en),
    .io_cfg_addr(gibs_42_io_cfg_addr),
    .io_cfg_data(gibs_42_io_cfg_data),
    .io_ipinNW_0(gibs_42_io_ipinNW_0),
    .io_ipinNW_1(gibs_42_io_ipinNW_1),
    .io_opinNW_0(gibs_42_io_opinNW_0),
    .io_ipinNE_0(gibs_42_io_ipinNE_0),
    .io_ipinNE_1(gibs_42_io_ipinNE_1),
    .io_opinNE_0(gibs_42_io_opinNE_0),
    .io_ipinSE_0(gibs_42_io_ipinSE_0),
    .io_ipinSE_1(gibs_42_io_ipinSE_1),
    .io_opinSE_0(gibs_42_io_opinSE_0),
    .io_ipinSW_0(gibs_42_io_ipinSW_0),
    .io_ipinSW_1(gibs_42_io_ipinSW_1),
    .io_opinSW_0(gibs_42_io_opinSW_0),
    .io_itrackW_0(gibs_42_io_itrackW_0),
    .io_otrackW_0(gibs_42_io_otrackW_0),
    .io_itrackN_0(gibs_42_io_itrackN_0),
    .io_otrackN_0(gibs_42_io_otrackN_0),
    .io_itrackE_0(gibs_42_io_itrackE_0),
    .io_otrackE_0(gibs_42_io_otrackE_0),
    .io_itrackS_0(gibs_42_io_itrackS_0),
    .io_otrackS_0(gibs_42_io_otrackS_0)
  );
  GIB_43 gibs_43 ( // @[CGRA.scala 333:21]
    .clock(gibs_43_clock),
    .reset(gibs_43_reset),
    .io_cfg_en(gibs_43_io_cfg_en),
    .io_cfg_addr(gibs_43_io_cfg_addr),
    .io_cfg_data(gibs_43_io_cfg_data),
    .io_ipinNW_0(gibs_43_io_ipinNW_0),
    .io_ipinNW_1(gibs_43_io_ipinNW_1),
    .io_opinNW_0(gibs_43_io_opinNW_0),
    .io_ipinNE_0(gibs_43_io_ipinNE_0),
    .io_opinNE_0(gibs_43_io_opinNE_0),
    .io_ipinSE_0(gibs_43_io_ipinSE_0),
    .io_opinSE_0(gibs_43_io_opinSE_0),
    .io_ipinSW_0(gibs_43_io_ipinSW_0),
    .io_ipinSW_1(gibs_43_io_ipinSW_1),
    .io_opinSW_0(gibs_43_io_opinSW_0),
    .io_itrackW_0(gibs_43_io_itrackW_0),
    .io_otrackW_0(gibs_43_io_otrackW_0),
    .io_itrackN_0(gibs_43_io_itrackN_0),
    .io_otrackN_0(gibs_43_io_otrackN_0),
    .io_itrackS_0(gibs_43_io_itrackS_0),
    .io_otrackS_0(gibs_43_io_otrackS_0)
  );
  GIB_44 gibs_44 ( // @[CGRA.scala 333:21]
    .clock(gibs_44_clock),
    .reset(gibs_44_reset),
    .io_cfg_en(gibs_44_io_cfg_en),
    .io_cfg_addr(gibs_44_io_cfg_addr),
    .io_cfg_data(gibs_44_io_cfg_data),
    .io_ipinNW_0(gibs_44_io_ipinNW_0),
    .io_opinNW_0(gibs_44_io_opinNW_0),
    .io_ipinNE_0(gibs_44_io_ipinNE_0),
    .io_ipinNE_1(gibs_44_io_ipinNE_1),
    .io_opinNE_0(gibs_44_io_opinNE_0),
    .io_ipinSE_0(gibs_44_io_ipinSE_0),
    .io_ipinSE_1(gibs_44_io_ipinSE_1),
    .io_opinSE_0(gibs_44_io_opinSE_0),
    .io_ipinSW_0(gibs_44_io_ipinSW_0),
    .io_opinSW_0(gibs_44_io_opinSW_0),
    .io_itrackN_0(gibs_44_io_itrackN_0),
    .io_otrackN_0(gibs_44_io_otrackN_0),
    .io_itrackE_0(gibs_44_io_itrackE_0),
    .io_otrackE_0(gibs_44_io_otrackE_0),
    .io_itrackS_0(gibs_44_io_itrackS_0),
    .io_otrackS_0(gibs_44_io_otrackS_0)
  );
  GIB_45 gibs_45 ( // @[CGRA.scala 333:21]
    .clock(gibs_45_clock),
    .reset(gibs_45_reset),
    .io_cfg_en(gibs_45_io_cfg_en),
    .io_cfg_addr(gibs_45_io_cfg_addr),
    .io_cfg_data(gibs_45_io_cfg_data),
    .io_ipinNW_0(gibs_45_io_ipinNW_0),
    .io_ipinNW_1(gibs_45_io_ipinNW_1),
    .io_opinNW_0(gibs_45_io_opinNW_0),
    .io_ipinNE_0(gibs_45_io_ipinNE_0),
    .io_ipinNE_1(gibs_45_io_ipinNE_1),
    .io_opinNE_0(gibs_45_io_opinNE_0),
    .io_ipinSE_0(gibs_45_io_ipinSE_0),
    .io_ipinSE_1(gibs_45_io_ipinSE_1),
    .io_opinSE_0(gibs_45_io_opinSE_0),
    .io_ipinSW_0(gibs_45_io_ipinSW_0),
    .io_ipinSW_1(gibs_45_io_ipinSW_1),
    .io_opinSW_0(gibs_45_io_opinSW_0),
    .io_itrackW_0(gibs_45_io_itrackW_0),
    .io_otrackW_0(gibs_45_io_otrackW_0),
    .io_itrackN_0(gibs_45_io_itrackN_0),
    .io_otrackN_0(gibs_45_io_otrackN_0),
    .io_itrackE_0(gibs_45_io_itrackE_0),
    .io_otrackE_0(gibs_45_io_otrackE_0),
    .io_itrackS_0(gibs_45_io_itrackS_0),
    .io_otrackS_0(gibs_45_io_otrackS_0)
  );
  GIB_46 gibs_46 ( // @[CGRA.scala 333:21]
    .clock(gibs_46_clock),
    .reset(gibs_46_reset),
    .io_cfg_en(gibs_46_io_cfg_en),
    .io_cfg_addr(gibs_46_io_cfg_addr),
    .io_cfg_data(gibs_46_io_cfg_data),
    .io_ipinNW_0(gibs_46_io_ipinNW_0),
    .io_ipinNW_1(gibs_46_io_ipinNW_1),
    .io_opinNW_0(gibs_46_io_opinNW_0),
    .io_ipinNE_0(gibs_46_io_ipinNE_0),
    .io_ipinNE_1(gibs_46_io_ipinNE_1),
    .io_opinNE_0(gibs_46_io_opinNE_0),
    .io_ipinSE_0(gibs_46_io_ipinSE_0),
    .io_ipinSE_1(gibs_46_io_ipinSE_1),
    .io_opinSE_0(gibs_46_io_opinSE_0),
    .io_ipinSW_0(gibs_46_io_ipinSW_0),
    .io_ipinSW_1(gibs_46_io_ipinSW_1),
    .io_opinSW_0(gibs_46_io_opinSW_0),
    .io_itrackW_0(gibs_46_io_itrackW_0),
    .io_otrackW_0(gibs_46_io_otrackW_0),
    .io_itrackN_0(gibs_46_io_itrackN_0),
    .io_otrackN_0(gibs_46_io_otrackN_0),
    .io_itrackE_0(gibs_46_io_itrackE_0),
    .io_otrackE_0(gibs_46_io_otrackE_0),
    .io_itrackS_0(gibs_46_io_itrackS_0),
    .io_otrackS_0(gibs_46_io_otrackS_0)
  );
  GIB_47 gibs_47 ( // @[CGRA.scala 333:21]
    .clock(gibs_47_clock),
    .reset(gibs_47_reset),
    .io_cfg_en(gibs_47_io_cfg_en),
    .io_cfg_addr(gibs_47_io_cfg_addr),
    .io_cfg_data(gibs_47_io_cfg_data),
    .io_ipinNW_0(gibs_47_io_ipinNW_0),
    .io_ipinNW_1(gibs_47_io_ipinNW_1),
    .io_opinNW_0(gibs_47_io_opinNW_0),
    .io_ipinNE_0(gibs_47_io_ipinNE_0),
    .io_opinNE_0(gibs_47_io_opinNE_0),
    .io_ipinSE_0(gibs_47_io_ipinSE_0),
    .io_opinSE_0(gibs_47_io_opinSE_0),
    .io_ipinSW_0(gibs_47_io_ipinSW_0),
    .io_ipinSW_1(gibs_47_io_ipinSW_1),
    .io_opinSW_0(gibs_47_io_opinSW_0),
    .io_itrackW_0(gibs_47_io_itrackW_0),
    .io_otrackW_0(gibs_47_io_otrackW_0),
    .io_itrackN_0(gibs_47_io_itrackN_0),
    .io_otrackN_0(gibs_47_io_otrackN_0),
    .io_itrackS_0(gibs_47_io_itrackS_0),
    .io_otrackS_0(gibs_47_io_otrackS_0)
  );
  GIB_48 gibs_48 ( // @[CGRA.scala 333:21]
    .clock(gibs_48_clock),
    .reset(gibs_48_reset),
    .io_cfg_en(gibs_48_io_cfg_en),
    .io_cfg_addr(gibs_48_io_cfg_addr),
    .io_cfg_data(gibs_48_io_cfg_data),
    .io_ipinNW_0(gibs_48_io_ipinNW_0),
    .io_opinNW_0(gibs_48_io_opinNW_0),
    .io_ipinNE_0(gibs_48_io_ipinNE_0),
    .io_ipinNE_1(gibs_48_io_ipinNE_1),
    .io_opinNE_0(gibs_48_io_opinNE_0),
    .io_ipinSE_0(gibs_48_io_ipinSE_0),
    .io_ipinSE_1(gibs_48_io_ipinSE_1),
    .io_opinSE_0(gibs_48_io_opinSE_0),
    .io_ipinSW_0(gibs_48_io_ipinSW_0),
    .io_opinSW_0(gibs_48_io_opinSW_0),
    .io_itrackN_0(gibs_48_io_itrackN_0),
    .io_otrackN_0(gibs_48_io_otrackN_0),
    .io_itrackE_0(gibs_48_io_itrackE_0),
    .io_otrackE_0(gibs_48_io_otrackE_0),
    .io_itrackS_0(gibs_48_io_itrackS_0),
    .io_otrackS_0(gibs_48_io_otrackS_0)
  );
  GIB_49 gibs_49 ( // @[CGRA.scala 333:21]
    .clock(gibs_49_clock),
    .reset(gibs_49_reset),
    .io_cfg_en(gibs_49_io_cfg_en),
    .io_cfg_addr(gibs_49_io_cfg_addr),
    .io_cfg_data(gibs_49_io_cfg_data),
    .io_ipinNW_0(gibs_49_io_ipinNW_0),
    .io_ipinNW_1(gibs_49_io_ipinNW_1),
    .io_opinNW_0(gibs_49_io_opinNW_0),
    .io_ipinNE_0(gibs_49_io_ipinNE_0),
    .io_ipinNE_1(gibs_49_io_ipinNE_1),
    .io_opinNE_0(gibs_49_io_opinNE_0),
    .io_ipinSE_0(gibs_49_io_ipinSE_0),
    .io_ipinSE_1(gibs_49_io_ipinSE_1),
    .io_opinSE_0(gibs_49_io_opinSE_0),
    .io_ipinSW_0(gibs_49_io_ipinSW_0),
    .io_ipinSW_1(gibs_49_io_ipinSW_1),
    .io_opinSW_0(gibs_49_io_opinSW_0),
    .io_itrackW_0(gibs_49_io_itrackW_0),
    .io_otrackW_0(gibs_49_io_otrackW_0),
    .io_itrackN_0(gibs_49_io_itrackN_0),
    .io_otrackN_0(gibs_49_io_otrackN_0),
    .io_itrackE_0(gibs_49_io_itrackE_0),
    .io_otrackE_0(gibs_49_io_otrackE_0),
    .io_itrackS_0(gibs_49_io_itrackS_0),
    .io_otrackS_0(gibs_49_io_otrackS_0)
  );
  GIB_50 gibs_50 ( // @[CGRA.scala 333:21]
    .clock(gibs_50_clock),
    .reset(gibs_50_reset),
    .io_cfg_en(gibs_50_io_cfg_en),
    .io_cfg_addr(gibs_50_io_cfg_addr),
    .io_cfg_data(gibs_50_io_cfg_data),
    .io_ipinNW_0(gibs_50_io_ipinNW_0),
    .io_ipinNW_1(gibs_50_io_ipinNW_1),
    .io_opinNW_0(gibs_50_io_opinNW_0),
    .io_ipinNE_0(gibs_50_io_ipinNE_0),
    .io_ipinNE_1(gibs_50_io_ipinNE_1),
    .io_opinNE_0(gibs_50_io_opinNE_0),
    .io_ipinSE_0(gibs_50_io_ipinSE_0),
    .io_ipinSE_1(gibs_50_io_ipinSE_1),
    .io_opinSE_0(gibs_50_io_opinSE_0),
    .io_ipinSW_0(gibs_50_io_ipinSW_0),
    .io_ipinSW_1(gibs_50_io_ipinSW_1),
    .io_opinSW_0(gibs_50_io_opinSW_0),
    .io_itrackW_0(gibs_50_io_itrackW_0),
    .io_otrackW_0(gibs_50_io_otrackW_0),
    .io_itrackN_0(gibs_50_io_itrackN_0),
    .io_otrackN_0(gibs_50_io_otrackN_0),
    .io_itrackE_0(gibs_50_io_itrackE_0),
    .io_otrackE_0(gibs_50_io_otrackE_0),
    .io_itrackS_0(gibs_50_io_itrackS_0),
    .io_otrackS_0(gibs_50_io_otrackS_0)
  );
  GIB_51 gibs_51 ( // @[CGRA.scala 333:21]
    .clock(gibs_51_clock),
    .reset(gibs_51_reset),
    .io_cfg_en(gibs_51_io_cfg_en),
    .io_cfg_addr(gibs_51_io_cfg_addr),
    .io_cfg_data(gibs_51_io_cfg_data),
    .io_ipinNW_0(gibs_51_io_ipinNW_0),
    .io_ipinNW_1(gibs_51_io_ipinNW_1),
    .io_opinNW_0(gibs_51_io_opinNW_0),
    .io_ipinNE_0(gibs_51_io_ipinNE_0),
    .io_opinNE_0(gibs_51_io_opinNE_0),
    .io_ipinSE_0(gibs_51_io_ipinSE_0),
    .io_opinSE_0(gibs_51_io_opinSE_0),
    .io_ipinSW_0(gibs_51_io_ipinSW_0),
    .io_ipinSW_1(gibs_51_io_ipinSW_1),
    .io_opinSW_0(gibs_51_io_opinSW_0),
    .io_itrackW_0(gibs_51_io_itrackW_0),
    .io_otrackW_0(gibs_51_io_otrackW_0),
    .io_itrackN_0(gibs_51_io_itrackN_0),
    .io_otrackN_0(gibs_51_io_otrackN_0),
    .io_itrackS_0(gibs_51_io_itrackS_0),
    .io_otrackS_0(gibs_51_io_otrackS_0)
  );
  GIB_52 gibs_52 ( // @[CGRA.scala 333:21]
    .clock(gibs_52_clock),
    .reset(gibs_52_reset),
    .io_cfg_en(gibs_52_io_cfg_en),
    .io_cfg_addr(gibs_52_io_cfg_addr),
    .io_cfg_data(gibs_52_io_cfg_data),
    .io_ipinNW_0(gibs_52_io_ipinNW_0),
    .io_opinNW_0(gibs_52_io_opinNW_0),
    .io_ipinNE_0(gibs_52_io_ipinNE_0),
    .io_ipinNE_1(gibs_52_io_ipinNE_1),
    .io_opinNE_0(gibs_52_io_opinNE_0),
    .io_ipinSE_0(gibs_52_io_ipinSE_0),
    .io_ipinSE_1(gibs_52_io_ipinSE_1),
    .io_opinSE_0(gibs_52_io_opinSE_0),
    .io_ipinSW_0(gibs_52_io_ipinSW_0),
    .io_opinSW_0(gibs_52_io_opinSW_0),
    .io_itrackN_0(gibs_52_io_itrackN_0),
    .io_otrackN_0(gibs_52_io_otrackN_0),
    .io_itrackE_0(gibs_52_io_itrackE_0),
    .io_otrackE_0(gibs_52_io_otrackE_0),
    .io_itrackS_0(gibs_52_io_itrackS_0),
    .io_otrackS_0(gibs_52_io_otrackS_0)
  );
  GIB_53 gibs_53 ( // @[CGRA.scala 333:21]
    .clock(gibs_53_clock),
    .reset(gibs_53_reset),
    .io_cfg_en(gibs_53_io_cfg_en),
    .io_cfg_addr(gibs_53_io_cfg_addr),
    .io_cfg_data(gibs_53_io_cfg_data),
    .io_ipinNW_0(gibs_53_io_ipinNW_0),
    .io_ipinNW_1(gibs_53_io_ipinNW_1),
    .io_opinNW_0(gibs_53_io_opinNW_0),
    .io_ipinNE_0(gibs_53_io_ipinNE_0),
    .io_ipinNE_1(gibs_53_io_ipinNE_1),
    .io_opinNE_0(gibs_53_io_opinNE_0),
    .io_ipinSE_0(gibs_53_io_ipinSE_0),
    .io_ipinSE_1(gibs_53_io_ipinSE_1),
    .io_opinSE_0(gibs_53_io_opinSE_0),
    .io_ipinSW_0(gibs_53_io_ipinSW_0),
    .io_ipinSW_1(gibs_53_io_ipinSW_1),
    .io_opinSW_0(gibs_53_io_opinSW_0),
    .io_itrackW_0(gibs_53_io_itrackW_0),
    .io_otrackW_0(gibs_53_io_otrackW_0),
    .io_itrackN_0(gibs_53_io_itrackN_0),
    .io_otrackN_0(gibs_53_io_otrackN_0),
    .io_itrackE_0(gibs_53_io_itrackE_0),
    .io_otrackE_0(gibs_53_io_otrackE_0),
    .io_itrackS_0(gibs_53_io_itrackS_0),
    .io_otrackS_0(gibs_53_io_otrackS_0)
  );
  GIB_54 gibs_54 ( // @[CGRA.scala 333:21]
    .clock(gibs_54_clock),
    .reset(gibs_54_reset),
    .io_cfg_en(gibs_54_io_cfg_en),
    .io_cfg_addr(gibs_54_io_cfg_addr),
    .io_cfg_data(gibs_54_io_cfg_data),
    .io_ipinNW_0(gibs_54_io_ipinNW_0),
    .io_ipinNW_1(gibs_54_io_ipinNW_1),
    .io_opinNW_0(gibs_54_io_opinNW_0),
    .io_ipinNE_0(gibs_54_io_ipinNE_0),
    .io_ipinNE_1(gibs_54_io_ipinNE_1),
    .io_opinNE_0(gibs_54_io_opinNE_0),
    .io_ipinSE_0(gibs_54_io_ipinSE_0),
    .io_ipinSE_1(gibs_54_io_ipinSE_1),
    .io_opinSE_0(gibs_54_io_opinSE_0),
    .io_ipinSW_0(gibs_54_io_ipinSW_0),
    .io_ipinSW_1(gibs_54_io_ipinSW_1),
    .io_opinSW_0(gibs_54_io_opinSW_0),
    .io_itrackW_0(gibs_54_io_itrackW_0),
    .io_otrackW_0(gibs_54_io_otrackW_0),
    .io_itrackN_0(gibs_54_io_itrackN_0),
    .io_otrackN_0(gibs_54_io_otrackN_0),
    .io_itrackE_0(gibs_54_io_itrackE_0),
    .io_otrackE_0(gibs_54_io_otrackE_0),
    .io_itrackS_0(gibs_54_io_itrackS_0),
    .io_otrackS_0(gibs_54_io_otrackS_0)
  );
  GIB_55 gibs_55 ( // @[CGRA.scala 333:21]
    .clock(gibs_55_clock),
    .reset(gibs_55_reset),
    .io_cfg_en(gibs_55_io_cfg_en),
    .io_cfg_addr(gibs_55_io_cfg_addr),
    .io_cfg_data(gibs_55_io_cfg_data),
    .io_ipinNW_0(gibs_55_io_ipinNW_0),
    .io_ipinNW_1(gibs_55_io_ipinNW_1),
    .io_opinNW_0(gibs_55_io_opinNW_0),
    .io_ipinNE_0(gibs_55_io_ipinNE_0),
    .io_opinNE_0(gibs_55_io_opinNE_0),
    .io_ipinSE_0(gibs_55_io_ipinSE_0),
    .io_opinSE_0(gibs_55_io_opinSE_0),
    .io_ipinSW_0(gibs_55_io_ipinSW_0),
    .io_ipinSW_1(gibs_55_io_ipinSW_1),
    .io_opinSW_0(gibs_55_io_opinSW_0),
    .io_itrackW_0(gibs_55_io_itrackW_0),
    .io_otrackW_0(gibs_55_io_otrackW_0),
    .io_itrackN_0(gibs_55_io_itrackN_0),
    .io_otrackN_0(gibs_55_io_otrackN_0),
    .io_itrackS_0(gibs_55_io_itrackS_0),
    .io_otrackS_0(gibs_55_io_otrackS_0)
  );
  GIB_56 gibs_56 ( // @[CGRA.scala 333:21]
    .clock(gibs_56_clock),
    .reset(gibs_56_reset),
    .io_cfg_en(gibs_56_io_cfg_en),
    .io_cfg_addr(gibs_56_io_cfg_addr),
    .io_cfg_data(gibs_56_io_cfg_data),
    .io_ipinNW_0(gibs_56_io_ipinNW_0),
    .io_opinNW_0(gibs_56_io_opinNW_0),
    .io_ipinNE_0(gibs_56_io_ipinNE_0),
    .io_ipinNE_1(gibs_56_io_ipinNE_1),
    .io_opinNE_0(gibs_56_io_opinNE_0),
    .io_ipinSE_0(gibs_56_io_ipinSE_0),
    .io_ipinSE_1(gibs_56_io_ipinSE_1),
    .io_opinSE_0(gibs_56_io_opinSE_0),
    .io_ipinSW_0(gibs_56_io_ipinSW_0),
    .io_opinSW_0(gibs_56_io_opinSW_0),
    .io_itrackN_0(gibs_56_io_itrackN_0),
    .io_otrackN_0(gibs_56_io_otrackN_0),
    .io_itrackE_0(gibs_56_io_itrackE_0),
    .io_otrackE_0(gibs_56_io_otrackE_0),
    .io_itrackS_0(gibs_56_io_itrackS_0),
    .io_otrackS_0(gibs_56_io_otrackS_0)
  );
  GIB_57 gibs_57 ( // @[CGRA.scala 333:21]
    .clock(gibs_57_clock),
    .reset(gibs_57_reset),
    .io_cfg_en(gibs_57_io_cfg_en),
    .io_cfg_addr(gibs_57_io_cfg_addr),
    .io_cfg_data(gibs_57_io_cfg_data),
    .io_ipinNW_0(gibs_57_io_ipinNW_0),
    .io_ipinNW_1(gibs_57_io_ipinNW_1),
    .io_opinNW_0(gibs_57_io_opinNW_0),
    .io_ipinNE_0(gibs_57_io_ipinNE_0),
    .io_ipinNE_1(gibs_57_io_ipinNE_1),
    .io_opinNE_0(gibs_57_io_opinNE_0),
    .io_ipinSE_0(gibs_57_io_ipinSE_0),
    .io_ipinSE_1(gibs_57_io_ipinSE_1),
    .io_opinSE_0(gibs_57_io_opinSE_0),
    .io_ipinSW_0(gibs_57_io_ipinSW_0),
    .io_ipinSW_1(gibs_57_io_ipinSW_1),
    .io_opinSW_0(gibs_57_io_opinSW_0),
    .io_itrackW_0(gibs_57_io_itrackW_0),
    .io_otrackW_0(gibs_57_io_otrackW_0),
    .io_itrackN_0(gibs_57_io_itrackN_0),
    .io_otrackN_0(gibs_57_io_otrackN_0),
    .io_itrackE_0(gibs_57_io_itrackE_0),
    .io_otrackE_0(gibs_57_io_otrackE_0),
    .io_itrackS_0(gibs_57_io_itrackS_0),
    .io_otrackS_0(gibs_57_io_otrackS_0)
  );
  GIB_58 gibs_58 ( // @[CGRA.scala 333:21]
    .clock(gibs_58_clock),
    .reset(gibs_58_reset),
    .io_cfg_en(gibs_58_io_cfg_en),
    .io_cfg_addr(gibs_58_io_cfg_addr),
    .io_cfg_data(gibs_58_io_cfg_data),
    .io_ipinNW_0(gibs_58_io_ipinNW_0),
    .io_ipinNW_1(gibs_58_io_ipinNW_1),
    .io_opinNW_0(gibs_58_io_opinNW_0),
    .io_ipinNE_0(gibs_58_io_ipinNE_0),
    .io_ipinNE_1(gibs_58_io_ipinNE_1),
    .io_opinNE_0(gibs_58_io_opinNE_0),
    .io_ipinSE_0(gibs_58_io_ipinSE_0),
    .io_ipinSE_1(gibs_58_io_ipinSE_1),
    .io_opinSE_0(gibs_58_io_opinSE_0),
    .io_ipinSW_0(gibs_58_io_ipinSW_0),
    .io_ipinSW_1(gibs_58_io_ipinSW_1),
    .io_opinSW_0(gibs_58_io_opinSW_0),
    .io_itrackW_0(gibs_58_io_itrackW_0),
    .io_otrackW_0(gibs_58_io_otrackW_0),
    .io_itrackN_0(gibs_58_io_itrackN_0),
    .io_otrackN_0(gibs_58_io_otrackN_0),
    .io_itrackE_0(gibs_58_io_itrackE_0),
    .io_otrackE_0(gibs_58_io_otrackE_0),
    .io_itrackS_0(gibs_58_io_itrackS_0),
    .io_otrackS_0(gibs_58_io_otrackS_0)
  );
  GIB_59 gibs_59 ( // @[CGRA.scala 333:21]
    .clock(gibs_59_clock),
    .reset(gibs_59_reset),
    .io_cfg_en(gibs_59_io_cfg_en),
    .io_cfg_addr(gibs_59_io_cfg_addr),
    .io_cfg_data(gibs_59_io_cfg_data),
    .io_ipinNW_0(gibs_59_io_ipinNW_0),
    .io_ipinNW_1(gibs_59_io_ipinNW_1),
    .io_opinNW_0(gibs_59_io_opinNW_0),
    .io_ipinNE_0(gibs_59_io_ipinNE_0),
    .io_opinNE_0(gibs_59_io_opinNE_0),
    .io_ipinSE_0(gibs_59_io_ipinSE_0),
    .io_opinSE_0(gibs_59_io_opinSE_0),
    .io_ipinSW_0(gibs_59_io_ipinSW_0),
    .io_ipinSW_1(gibs_59_io_ipinSW_1),
    .io_opinSW_0(gibs_59_io_opinSW_0),
    .io_itrackW_0(gibs_59_io_itrackW_0),
    .io_otrackW_0(gibs_59_io_otrackW_0),
    .io_itrackN_0(gibs_59_io_itrackN_0),
    .io_otrackN_0(gibs_59_io_otrackN_0),
    .io_itrackS_0(gibs_59_io_itrackS_0),
    .io_otrackS_0(gibs_59_io_otrackS_0)
  );
  GIB_60 gibs_60 ( // @[CGRA.scala 333:21]
    .clock(gibs_60_clock),
    .reset(gibs_60_reset),
    .io_cfg_en(gibs_60_io_cfg_en),
    .io_cfg_addr(gibs_60_io_cfg_addr),
    .io_cfg_data(gibs_60_io_cfg_data),
    .io_ipinNW_0(gibs_60_io_ipinNW_0),
    .io_opinNW_0(gibs_60_io_opinNW_0),
    .io_ipinNE_0(gibs_60_io_ipinNE_0),
    .io_ipinNE_1(gibs_60_io_ipinNE_1),
    .io_opinNE_0(gibs_60_io_opinNE_0),
    .io_ipinSE_0(gibs_60_io_ipinSE_0),
    .io_ipinSE_1(gibs_60_io_ipinSE_1),
    .io_opinSE_0(gibs_60_io_opinSE_0),
    .io_ipinSW_0(gibs_60_io_ipinSW_0),
    .io_opinSW_0(gibs_60_io_opinSW_0),
    .io_itrackN_0(gibs_60_io_itrackN_0),
    .io_otrackN_0(gibs_60_io_otrackN_0),
    .io_itrackE_0(gibs_60_io_itrackE_0),
    .io_otrackE_0(gibs_60_io_otrackE_0),
    .io_itrackS_0(gibs_60_io_itrackS_0),
    .io_otrackS_0(gibs_60_io_otrackS_0)
  );
  GIB_61 gibs_61 ( // @[CGRA.scala 333:21]
    .clock(gibs_61_clock),
    .reset(gibs_61_reset),
    .io_cfg_en(gibs_61_io_cfg_en),
    .io_cfg_addr(gibs_61_io_cfg_addr),
    .io_cfg_data(gibs_61_io_cfg_data),
    .io_ipinNW_0(gibs_61_io_ipinNW_0),
    .io_ipinNW_1(gibs_61_io_ipinNW_1),
    .io_opinNW_0(gibs_61_io_opinNW_0),
    .io_ipinNE_0(gibs_61_io_ipinNE_0),
    .io_ipinNE_1(gibs_61_io_ipinNE_1),
    .io_opinNE_0(gibs_61_io_opinNE_0),
    .io_ipinSE_0(gibs_61_io_ipinSE_0),
    .io_ipinSE_1(gibs_61_io_ipinSE_1),
    .io_opinSE_0(gibs_61_io_opinSE_0),
    .io_ipinSW_0(gibs_61_io_ipinSW_0),
    .io_ipinSW_1(gibs_61_io_ipinSW_1),
    .io_opinSW_0(gibs_61_io_opinSW_0),
    .io_itrackW_0(gibs_61_io_itrackW_0),
    .io_otrackW_0(gibs_61_io_otrackW_0),
    .io_itrackN_0(gibs_61_io_itrackN_0),
    .io_otrackN_0(gibs_61_io_otrackN_0),
    .io_itrackE_0(gibs_61_io_itrackE_0),
    .io_otrackE_0(gibs_61_io_otrackE_0),
    .io_itrackS_0(gibs_61_io_itrackS_0),
    .io_otrackS_0(gibs_61_io_otrackS_0)
  );
  GIB_62 gibs_62 ( // @[CGRA.scala 333:21]
    .clock(gibs_62_clock),
    .reset(gibs_62_reset),
    .io_cfg_en(gibs_62_io_cfg_en),
    .io_cfg_addr(gibs_62_io_cfg_addr),
    .io_cfg_data(gibs_62_io_cfg_data),
    .io_ipinNW_0(gibs_62_io_ipinNW_0),
    .io_ipinNW_1(gibs_62_io_ipinNW_1),
    .io_opinNW_0(gibs_62_io_opinNW_0),
    .io_ipinNE_0(gibs_62_io_ipinNE_0),
    .io_ipinNE_1(gibs_62_io_ipinNE_1),
    .io_opinNE_0(gibs_62_io_opinNE_0),
    .io_ipinSE_0(gibs_62_io_ipinSE_0),
    .io_ipinSE_1(gibs_62_io_ipinSE_1),
    .io_opinSE_0(gibs_62_io_opinSE_0),
    .io_ipinSW_0(gibs_62_io_ipinSW_0),
    .io_ipinSW_1(gibs_62_io_ipinSW_1),
    .io_opinSW_0(gibs_62_io_opinSW_0),
    .io_itrackW_0(gibs_62_io_itrackW_0),
    .io_otrackW_0(gibs_62_io_otrackW_0),
    .io_itrackN_0(gibs_62_io_itrackN_0),
    .io_otrackN_0(gibs_62_io_otrackN_0),
    .io_itrackE_0(gibs_62_io_itrackE_0),
    .io_otrackE_0(gibs_62_io_otrackE_0),
    .io_itrackS_0(gibs_62_io_itrackS_0),
    .io_otrackS_0(gibs_62_io_otrackS_0)
  );
  GIB_63 gibs_63 ( // @[CGRA.scala 333:21]
    .clock(gibs_63_clock),
    .reset(gibs_63_reset),
    .io_cfg_en(gibs_63_io_cfg_en),
    .io_cfg_addr(gibs_63_io_cfg_addr),
    .io_cfg_data(gibs_63_io_cfg_data),
    .io_ipinNW_0(gibs_63_io_ipinNW_0),
    .io_ipinNW_1(gibs_63_io_ipinNW_1),
    .io_opinNW_0(gibs_63_io_opinNW_0),
    .io_ipinNE_0(gibs_63_io_ipinNE_0),
    .io_opinNE_0(gibs_63_io_opinNE_0),
    .io_ipinSE_0(gibs_63_io_ipinSE_0),
    .io_opinSE_0(gibs_63_io_opinSE_0),
    .io_ipinSW_0(gibs_63_io_ipinSW_0),
    .io_ipinSW_1(gibs_63_io_ipinSW_1),
    .io_opinSW_0(gibs_63_io_opinSW_0),
    .io_itrackW_0(gibs_63_io_itrackW_0),
    .io_otrackW_0(gibs_63_io_otrackW_0),
    .io_itrackN_0(gibs_63_io_itrackN_0),
    .io_otrackN_0(gibs_63_io_otrackN_0),
    .io_itrackS_0(gibs_63_io_itrackS_0),
    .io_otrackS_0(gibs_63_io_otrackS_0)
  );
  GIB_64 gibs_64 ( // @[CGRA.scala 333:21]
    .clock(gibs_64_clock),
    .reset(gibs_64_reset),
    .io_cfg_en(gibs_64_io_cfg_en),
    .io_cfg_addr(gibs_64_io_cfg_addr),
    .io_cfg_data(gibs_64_io_cfg_data),
    .io_ipinNW_0(gibs_64_io_ipinNW_0),
    .io_opinNW_0(gibs_64_io_opinNW_0),
    .io_ipinNE_0(gibs_64_io_ipinNE_0),
    .io_ipinNE_1(gibs_64_io_ipinNE_1),
    .io_opinNE_0(gibs_64_io_opinNE_0),
    .io_ipinSE_0(gibs_64_io_ipinSE_0),
    .io_ipinSE_1(gibs_64_io_ipinSE_1),
    .io_opinSE_0(gibs_64_io_opinSE_0),
    .io_ipinSW_0(gibs_64_io_ipinSW_0),
    .io_opinSW_0(gibs_64_io_opinSW_0),
    .io_itrackN_0(gibs_64_io_itrackN_0),
    .io_otrackN_0(gibs_64_io_otrackN_0),
    .io_itrackE_0(gibs_64_io_itrackE_0),
    .io_otrackE_0(gibs_64_io_otrackE_0),
    .io_itrackS_0(gibs_64_io_itrackS_0),
    .io_otrackS_0(gibs_64_io_otrackS_0)
  );
  GIB_65 gibs_65 ( // @[CGRA.scala 333:21]
    .clock(gibs_65_clock),
    .reset(gibs_65_reset),
    .io_cfg_en(gibs_65_io_cfg_en),
    .io_cfg_addr(gibs_65_io_cfg_addr),
    .io_cfg_data(gibs_65_io_cfg_data),
    .io_ipinNW_0(gibs_65_io_ipinNW_0),
    .io_ipinNW_1(gibs_65_io_ipinNW_1),
    .io_opinNW_0(gibs_65_io_opinNW_0),
    .io_ipinNE_0(gibs_65_io_ipinNE_0),
    .io_ipinNE_1(gibs_65_io_ipinNE_1),
    .io_opinNE_0(gibs_65_io_opinNE_0),
    .io_ipinSE_0(gibs_65_io_ipinSE_0),
    .io_ipinSE_1(gibs_65_io_ipinSE_1),
    .io_opinSE_0(gibs_65_io_opinSE_0),
    .io_ipinSW_0(gibs_65_io_ipinSW_0),
    .io_ipinSW_1(gibs_65_io_ipinSW_1),
    .io_opinSW_0(gibs_65_io_opinSW_0),
    .io_itrackW_0(gibs_65_io_itrackW_0),
    .io_otrackW_0(gibs_65_io_otrackW_0),
    .io_itrackN_0(gibs_65_io_itrackN_0),
    .io_otrackN_0(gibs_65_io_otrackN_0),
    .io_itrackE_0(gibs_65_io_itrackE_0),
    .io_otrackE_0(gibs_65_io_otrackE_0),
    .io_itrackS_0(gibs_65_io_itrackS_0),
    .io_otrackS_0(gibs_65_io_otrackS_0)
  );
  GIB_66 gibs_66 ( // @[CGRA.scala 333:21]
    .clock(gibs_66_clock),
    .reset(gibs_66_reset),
    .io_cfg_en(gibs_66_io_cfg_en),
    .io_cfg_addr(gibs_66_io_cfg_addr),
    .io_cfg_data(gibs_66_io_cfg_data),
    .io_ipinNW_0(gibs_66_io_ipinNW_0),
    .io_ipinNW_1(gibs_66_io_ipinNW_1),
    .io_opinNW_0(gibs_66_io_opinNW_0),
    .io_ipinNE_0(gibs_66_io_ipinNE_0),
    .io_ipinNE_1(gibs_66_io_ipinNE_1),
    .io_opinNE_0(gibs_66_io_opinNE_0),
    .io_ipinSE_0(gibs_66_io_ipinSE_0),
    .io_ipinSE_1(gibs_66_io_ipinSE_1),
    .io_opinSE_0(gibs_66_io_opinSE_0),
    .io_ipinSW_0(gibs_66_io_ipinSW_0),
    .io_ipinSW_1(gibs_66_io_ipinSW_1),
    .io_opinSW_0(gibs_66_io_opinSW_0),
    .io_itrackW_0(gibs_66_io_itrackW_0),
    .io_otrackW_0(gibs_66_io_otrackW_0),
    .io_itrackN_0(gibs_66_io_itrackN_0),
    .io_otrackN_0(gibs_66_io_otrackN_0),
    .io_itrackE_0(gibs_66_io_itrackE_0),
    .io_otrackE_0(gibs_66_io_otrackE_0),
    .io_itrackS_0(gibs_66_io_itrackS_0),
    .io_otrackS_0(gibs_66_io_otrackS_0)
  );
  GIB_67 gibs_67 ( // @[CGRA.scala 333:21]
    .clock(gibs_67_clock),
    .reset(gibs_67_reset),
    .io_cfg_en(gibs_67_io_cfg_en),
    .io_cfg_addr(gibs_67_io_cfg_addr),
    .io_cfg_data(gibs_67_io_cfg_data),
    .io_ipinNW_0(gibs_67_io_ipinNW_0),
    .io_ipinNW_1(gibs_67_io_ipinNW_1),
    .io_opinNW_0(gibs_67_io_opinNW_0),
    .io_ipinNE_0(gibs_67_io_ipinNE_0),
    .io_opinNE_0(gibs_67_io_opinNE_0),
    .io_ipinSE_0(gibs_67_io_ipinSE_0),
    .io_opinSE_0(gibs_67_io_opinSE_0),
    .io_ipinSW_0(gibs_67_io_ipinSW_0),
    .io_ipinSW_1(gibs_67_io_ipinSW_1),
    .io_opinSW_0(gibs_67_io_opinSW_0),
    .io_itrackW_0(gibs_67_io_itrackW_0),
    .io_otrackW_0(gibs_67_io_otrackW_0),
    .io_itrackN_0(gibs_67_io_itrackN_0),
    .io_otrackN_0(gibs_67_io_otrackN_0),
    .io_itrackS_0(gibs_67_io_itrackS_0),
    .io_otrackS_0(gibs_67_io_otrackS_0)
  );
  GIB_68 gibs_68 ( // @[CGRA.scala 333:21]
    .clock(gibs_68_clock),
    .reset(gibs_68_reset),
    .io_cfg_en(gibs_68_io_cfg_en),
    .io_cfg_addr(gibs_68_io_cfg_addr),
    .io_cfg_data(gibs_68_io_cfg_data),
    .io_ipinNW_0(gibs_68_io_ipinNW_0),
    .io_opinNW_0(gibs_68_io_opinNW_0),
    .io_ipinNE_0(gibs_68_io_ipinNE_0),
    .io_ipinNE_1(gibs_68_io_ipinNE_1),
    .io_opinNE_0(gibs_68_io_opinNE_0),
    .io_ipinSE_0(gibs_68_io_ipinSE_0),
    .io_ipinSE_1(gibs_68_io_ipinSE_1),
    .io_opinSE_0(gibs_68_io_opinSE_0),
    .io_ipinSW_0(gibs_68_io_ipinSW_0),
    .io_opinSW_0(gibs_68_io_opinSW_0),
    .io_itrackN_0(gibs_68_io_itrackN_0),
    .io_otrackN_0(gibs_68_io_otrackN_0),
    .io_itrackE_0(gibs_68_io_itrackE_0),
    .io_otrackE_0(gibs_68_io_otrackE_0),
    .io_itrackS_0(gibs_68_io_itrackS_0),
    .io_otrackS_0(gibs_68_io_otrackS_0)
  );
  GIB_69 gibs_69 ( // @[CGRA.scala 333:21]
    .clock(gibs_69_clock),
    .reset(gibs_69_reset),
    .io_cfg_en(gibs_69_io_cfg_en),
    .io_cfg_addr(gibs_69_io_cfg_addr),
    .io_cfg_data(gibs_69_io_cfg_data),
    .io_ipinNW_0(gibs_69_io_ipinNW_0),
    .io_ipinNW_1(gibs_69_io_ipinNW_1),
    .io_opinNW_0(gibs_69_io_opinNW_0),
    .io_ipinNE_0(gibs_69_io_ipinNE_0),
    .io_ipinNE_1(gibs_69_io_ipinNE_1),
    .io_opinNE_0(gibs_69_io_opinNE_0),
    .io_ipinSE_0(gibs_69_io_ipinSE_0),
    .io_ipinSE_1(gibs_69_io_ipinSE_1),
    .io_opinSE_0(gibs_69_io_opinSE_0),
    .io_ipinSW_0(gibs_69_io_ipinSW_0),
    .io_ipinSW_1(gibs_69_io_ipinSW_1),
    .io_opinSW_0(gibs_69_io_opinSW_0),
    .io_itrackW_0(gibs_69_io_itrackW_0),
    .io_otrackW_0(gibs_69_io_otrackW_0),
    .io_itrackN_0(gibs_69_io_itrackN_0),
    .io_otrackN_0(gibs_69_io_otrackN_0),
    .io_itrackE_0(gibs_69_io_itrackE_0),
    .io_otrackE_0(gibs_69_io_otrackE_0),
    .io_itrackS_0(gibs_69_io_itrackS_0),
    .io_otrackS_0(gibs_69_io_otrackS_0)
  );
  GIB_70 gibs_70 ( // @[CGRA.scala 333:21]
    .clock(gibs_70_clock),
    .reset(gibs_70_reset),
    .io_cfg_en(gibs_70_io_cfg_en),
    .io_cfg_addr(gibs_70_io_cfg_addr),
    .io_cfg_data(gibs_70_io_cfg_data),
    .io_ipinNW_0(gibs_70_io_ipinNW_0),
    .io_ipinNW_1(gibs_70_io_ipinNW_1),
    .io_opinNW_0(gibs_70_io_opinNW_0),
    .io_ipinNE_0(gibs_70_io_ipinNE_0),
    .io_ipinNE_1(gibs_70_io_ipinNE_1),
    .io_opinNE_0(gibs_70_io_opinNE_0),
    .io_ipinSE_0(gibs_70_io_ipinSE_0),
    .io_ipinSE_1(gibs_70_io_ipinSE_1),
    .io_opinSE_0(gibs_70_io_opinSE_0),
    .io_ipinSW_0(gibs_70_io_ipinSW_0),
    .io_ipinSW_1(gibs_70_io_ipinSW_1),
    .io_opinSW_0(gibs_70_io_opinSW_0),
    .io_itrackW_0(gibs_70_io_itrackW_0),
    .io_otrackW_0(gibs_70_io_otrackW_0),
    .io_itrackN_0(gibs_70_io_itrackN_0),
    .io_otrackN_0(gibs_70_io_otrackN_0),
    .io_itrackE_0(gibs_70_io_itrackE_0),
    .io_otrackE_0(gibs_70_io_otrackE_0),
    .io_itrackS_0(gibs_70_io_itrackS_0),
    .io_otrackS_0(gibs_70_io_otrackS_0)
  );
  GIB_71 gibs_71 ( // @[CGRA.scala 333:21]
    .clock(gibs_71_clock),
    .reset(gibs_71_reset),
    .io_cfg_en(gibs_71_io_cfg_en),
    .io_cfg_addr(gibs_71_io_cfg_addr),
    .io_cfg_data(gibs_71_io_cfg_data),
    .io_ipinNW_0(gibs_71_io_ipinNW_0),
    .io_ipinNW_1(gibs_71_io_ipinNW_1),
    .io_opinNW_0(gibs_71_io_opinNW_0),
    .io_ipinNE_0(gibs_71_io_ipinNE_0),
    .io_opinNE_0(gibs_71_io_opinNE_0),
    .io_ipinSE_0(gibs_71_io_ipinSE_0),
    .io_opinSE_0(gibs_71_io_opinSE_0),
    .io_ipinSW_0(gibs_71_io_ipinSW_0),
    .io_ipinSW_1(gibs_71_io_ipinSW_1),
    .io_opinSW_0(gibs_71_io_opinSW_0),
    .io_itrackW_0(gibs_71_io_itrackW_0),
    .io_otrackW_0(gibs_71_io_otrackW_0),
    .io_itrackN_0(gibs_71_io_itrackN_0),
    .io_otrackN_0(gibs_71_io_otrackN_0),
    .io_itrackS_0(gibs_71_io_itrackS_0),
    .io_otrackS_0(gibs_71_io_otrackS_0)
  );
  GIB_72 gibs_72 ( // @[CGRA.scala 333:21]
    .clock(gibs_72_clock),
    .reset(gibs_72_reset),
    .io_cfg_en(gibs_72_io_cfg_en),
    .io_cfg_addr(gibs_72_io_cfg_addr),
    .io_cfg_data(gibs_72_io_cfg_data),
    .io_ipinNW_0(gibs_72_io_ipinNW_0),
    .io_opinNW_0(gibs_72_io_opinNW_0),
    .io_ipinNE_0(gibs_72_io_ipinNE_0),
    .io_ipinNE_1(gibs_72_io_ipinNE_1),
    .io_opinNE_0(gibs_72_io_opinNE_0),
    .io_ipinSE_0(gibs_72_io_ipinSE_0),
    .io_ipinSE_1(gibs_72_io_ipinSE_1),
    .io_opinSE_0(gibs_72_io_opinSE_0),
    .io_ipinSW_0(gibs_72_io_ipinSW_0),
    .io_opinSW_0(gibs_72_io_opinSW_0),
    .io_itrackN_0(gibs_72_io_itrackN_0),
    .io_otrackN_0(gibs_72_io_otrackN_0),
    .io_itrackE_0(gibs_72_io_itrackE_0),
    .io_otrackE_0(gibs_72_io_otrackE_0),
    .io_itrackS_0(gibs_72_io_itrackS_0),
    .io_otrackS_0(gibs_72_io_otrackS_0)
  );
  GIB_73 gibs_73 ( // @[CGRA.scala 333:21]
    .clock(gibs_73_clock),
    .reset(gibs_73_reset),
    .io_cfg_en(gibs_73_io_cfg_en),
    .io_cfg_addr(gibs_73_io_cfg_addr),
    .io_cfg_data(gibs_73_io_cfg_data),
    .io_ipinNW_0(gibs_73_io_ipinNW_0),
    .io_ipinNW_1(gibs_73_io_ipinNW_1),
    .io_opinNW_0(gibs_73_io_opinNW_0),
    .io_ipinNE_0(gibs_73_io_ipinNE_0),
    .io_ipinNE_1(gibs_73_io_ipinNE_1),
    .io_opinNE_0(gibs_73_io_opinNE_0),
    .io_ipinSE_0(gibs_73_io_ipinSE_0),
    .io_ipinSE_1(gibs_73_io_ipinSE_1),
    .io_opinSE_0(gibs_73_io_opinSE_0),
    .io_ipinSW_0(gibs_73_io_ipinSW_0),
    .io_ipinSW_1(gibs_73_io_ipinSW_1),
    .io_opinSW_0(gibs_73_io_opinSW_0),
    .io_itrackW_0(gibs_73_io_itrackW_0),
    .io_otrackW_0(gibs_73_io_otrackW_0),
    .io_itrackN_0(gibs_73_io_itrackN_0),
    .io_otrackN_0(gibs_73_io_otrackN_0),
    .io_itrackE_0(gibs_73_io_itrackE_0),
    .io_otrackE_0(gibs_73_io_otrackE_0),
    .io_itrackS_0(gibs_73_io_itrackS_0),
    .io_otrackS_0(gibs_73_io_otrackS_0)
  );
  GIB_74 gibs_74 ( // @[CGRA.scala 333:21]
    .clock(gibs_74_clock),
    .reset(gibs_74_reset),
    .io_cfg_en(gibs_74_io_cfg_en),
    .io_cfg_addr(gibs_74_io_cfg_addr),
    .io_cfg_data(gibs_74_io_cfg_data),
    .io_ipinNW_0(gibs_74_io_ipinNW_0),
    .io_ipinNW_1(gibs_74_io_ipinNW_1),
    .io_opinNW_0(gibs_74_io_opinNW_0),
    .io_ipinNE_0(gibs_74_io_ipinNE_0),
    .io_ipinNE_1(gibs_74_io_ipinNE_1),
    .io_opinNE_0(gibs_74_io_opinNE_0),
    .io_ipinSE_0(gibs_74_io_ipinSE_0),
    .io_ipinSE_1(gibs_74_io_ipinSE_1),
    .io_opinSE_0(gibs_74_io_opinSE_0),
    .io_ipinSW_0(gibs_74_io_ipinSW_0),
    .io_ipinSW_1(gibs_74_io_ipinSW_1),
    .io_opinSW_0(gibs_74_io_opinSW_0),
    .io_itrackW_0(gibs_74_io_itrackW_0),
    .io_otrackW_0(gibs_74_io_otrackW_0),
    .io_itrackN_0(gibs_74_io_itrackN_0),
    .io_otrackN_0(gibs_74_io_otrackN_0),
    .io_itrackE_0(gibs_74_io_itrackE_0),
    .io_otrackE_0(gibs_74_io_otrackE_0),
    .io_itrackS_0(gibs_74_io_itrackS_0),
    .io_otrackS_0(gibs_74_io_otrackS_0)
  );
  GIB_75 gibs_75 ( // @[CGRA.scala 333:21]
    .clock(gibs_75_clock),
    .reset(gibs_75_reset),
    .io_cfg_en(gibs_75_io_cfg_en),
    .io_cfg_addr(gibs_75_io_cfg_addr),
    .io_cfg_data(gibs_75_io_cfg_data),
    .io_ipinNW_0(gibs_75_io_ipinNW_0),
    .io_ipinNW_1(gibs_75_io_ipinNW_1),
    .io_opinNW_0(gibs_75_io_opinNW_0),
    .io_ipinNE_0(gibs_75_io_ipinNE_0),
    .io_opinNE_0(gibs_75_io_opinNE_0),
    .io_ipinSE_0(gibs_75_io_ipinSE_0),
    .io_opinSE_0(gibs_75_io_opinSE_0),
    .io_ipinSW_0(gibs_75_io_ipinSW_0),
    .io_ipinSW_1(gibs_75_io_ipinSW_1),
    .io_opinSW_0(gibs_75_io_opinSW_0),
    .io_itrackW_0(gibs_75_io_itrackW_0),
    .io_otrackW_0(gibs_75_io_otrackW_0),
    .io_itrackN_0(gibs_75_io_itrackN_0),
    .io_otrackN_0(gibs_75_io_otrackN_0),
    .io_itrackS_0(gibs_75_io_itrackS_0),
    .io_otrackS_0(gibs_75_io_otrackS_0)
  );
  GIB_76 gibs_76 ( // @[CGRA.scala 333:21]
    .clock(gibs_76_clock),
    .reset(gibs_76_reset),
    .io_cfg_en(gibs_76_io_cfg_en),
    .io_cfg_addr(gibs_76_io_cfg_addr),
    .io_cfg_data(gibs_76_io_cfg_data),
    .io_ipinNW_0(gibs_76_io_ipinNW_0),
    .io_opinNW_0(gibs_76_io_opinNW_0),
    .io_ipinNE_0(gibs_76_io_ipinNE_0),
    .io_ipinNE_1(gibs_76_io_ipinNE_1),
    .io_opinNE_0(gibs_76_io_opinNE_0),
    .io_ipinSE_0(gibs_76_io_ipinSE_0),
    .io_opinSE_0(gibs_76_io_opinSE_0),
    .io_itrackN_0(gibs_76_io_itrackN_0),
    .io_otrackN_0(gibs_76_io_otrackN_0),
    .io_itrackE_0(gibs_76_io_itrackE_0),
    .io_otrackE_0(gibs_76_io_otrackE_0)
  );
  GIB_77 gibs_77 ( // @[CGRA.scala 333:21]
    .clock(gibs_77_clock),
    .reset(gibs_77_reset),
    .io_cfg_en(gibs_77_io_cfg_en),
    .io_cfg_addr(gibs_77_io_cfg_addr),
    .io_cfg_data(gibs_77_io_cfg_data),
    .io_ipinNW_0(gibs_77_io_ipinNW_0),
    .io_ipinNW_1(gibs_77_io_ipinNW_1),
    .io_opinNW_0(gibs_77_io_opinNW_0),
    .io_ipinNE_0(gibs_77_io_ipinNE_0),
    .io_ipinNE_1(gibs_77_io_ipinNE_1),
    .io_opinNE_0(gibs_77_io_opinNE_0),
    .io_ipinSE_0(gibs_77_io_ipinSE_0),
    .io_opinSE_0(gibs_77_io_opinSE_0),
    .io_ipinSW_0(gibs_77_io_ipinSW_0),
    .io_opinSW_0(gibs_77_io_opinSW_0),
    .io_itrackW_0(gibs_77_io_itrackW_0),
    .io_otrackW_0(gibs_77_io_otrackW_0),
    .io_itrackN_0(gibs_77_io_itrackN_0),
    .io_otrackN_0(gibs_77_io_otrackN_0),
    .io_itrackE_0(gibs_77_io_itrackE_0),
    .io_otrackE_0(gibs_77_io_otrackE_0)
  );
  GIB_78 gibs_78 ( // @[CGRA.scala 333:21]
    .clock(gibs_78_clock),
    .reset(gibs_78_reset),
    .io_cfg_en(gibs_78_io_cfg_en),
    .io_cfg_addr(gibs_78_io_cfg_addr),
    .io_cfg_data(gibs_78_io_cfg_data),
    .io_ipinNW_0(gibs_78_io_ipinNW_0),
    .io_ipinNW_1(gibs_78_io_ipinNW_1),
    .io_opinNW_0(gibs_78_io_opinNW_0),
    .io_ipinNE_0(gibs_78_io_ipinNE_0),
    .io_ipinNE_1(gibs_78_io_ipinNE_1),
    .io_opinNE_0(gibs_78_io_opinNE_0),
    .io_ipinSE_0(gibs_78_io_ipinSE_0),
    .io_opinSE_0(gibs_78_io_opinSE_0),
    .io_ipinSW_0(gibs_78_io_ipinSW_0),
    .io_opinSW_0(gibs_78_io_opinSW_0),
    .io_itrackW_0(gibs_78_io_itrackW_0),
    .io_otrackW_0(gibs_78_io_otrackW_0),
    .io_itrackN_0(gibs_78_io_itrackN_0),
    .io_otrackN_0(gibs_78_io_otrackN_0),
    .io_itrackE_0(gibs_78_io_itrackE_0),
    .io_otrackE_0(gibs_78_io_otrackE_0)
  );
  GIB_79 gibs_79 ( // @[CGRA.scala 333:21]
    .clock(gibs_79_clock),
    .reset(gibs_79_reset),
    .io_cfg_en(gibs_79_io_cfg_en),
    .io_cfg_addr(gibs_79_io_cfg_addr),
    .io_cfg_data(gibs_79_io_cfg_data),
    .io_ipinNW_0(gibs_79_io_ipinNW_0),
    .io_ipinNW_1(gibs_79_io_ipinNW_1),
    .io_opinNW_0(gibs_79_io_opinNW_0),
    .io_ipinNE_0(gibs_79_io_ipinNE_0),
    .io_opinNE_0(gibs_79_io_opinNE_0),
    .io_ipinSW_0(gibs_79_io_ipinSW_0),
    .io_opinSW_0(gibs_79_io_opinSW_0),
    .io_itrackW_0(gibs_79_io_itrackW_0),
    .io_otrackW_0(gibs_79_io_otrackW_0),
    .io_itrackN_0(gibs_79_io_itrackN_0),
    .io_otrackN_0(gibs_79_io_otrackN_0)
  );
  LSU lsus_0 ( // @[CGRA.scala 364:21]
    .clock(lsus_0_clock),
    .reset(lsus_0_reset),
    .io_cfg_en(lsus_0_io_cfg_en),
    .io_cfg_addr(lsus_0_io_cfg_addr),
    .io_cfg_data(lsus_0_io_cfg_data),
    .io_hostInterface_read_addr(lsus_0_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_0_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_0_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_0_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_0_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_0_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_0_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_0_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_0_io_hostInterface_cycle),
    .io_en(lsus_0_io_en),
    .io_in_0(lsus_0_io_in_0),
    .io_in_1(lsus_0_io_in_1),
    .io_out_0(lsus_0_io_out_0)
  );
  LSU_1 lsus_1 ( // @[CGRA.scala 364:21]
    .clock(lsus_1_clock),
    .reset(lsus_1_reset),
    .io_cfg_en(lsus_1_io_cfg_en),
    .io_cfg_addr(lsus_1_io_cfg_addr),
    .io_cfg_data(lsus_1_io_cfg_data),
    .io_hostInterface_read_addr(lsus_1_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_1_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_1_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_1_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_1_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_1_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_1_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_1_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_1_io_hostInterface_cycle),
    .io_en(lsus_1_io_en),
    .io_in_0(lsus_1_io_in_0),
    .io_in_1(lsus_1_io_in_1),
    .io_out_0(lsus_1_io_out_0)
  );
  LSU_2 lsus_2 ( // @[CGRA.scala 364:21]
    .clock(lsus_2_clock),
    .reset(lsus_2_reset),
    .io_cfg_en(lsus_2_io_cfg_en),
    .io_cfg_addr(lsus_2_io_cfg_addr),
    .io_cfg_data(lsus_2_io_cfg_data),
    .io_hostInterface_read_addr(lsus_2_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_2_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_2_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_2_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_2_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_2_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_2_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_2_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_2_io_hostInterface_cycle),
    .io_en(lsus_2_io_en),
    .io_in_0(lsus_2_io_in_0),
    .io_in_1(lsus_2_io_in_1),
    .io_out_0(lsus_2_io_out_0)
  );
  LSU_3 lsus_3 ( // @[CGRA.scala 364:21]
    .clock(lsus_3_clock),
    .reset(lsus_3_reset),
    .io_cfg_en(lsus_3_io_cfg_en),
    .io_cfg_addr(lsus_3_io_cfg_addr),
    .io_cfg_data(lsus_3_io_cfg_data),
    .io_hostInterface_read_addr(lsus_3_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_3_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_3_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_3_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_3_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_3_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_3_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_3_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_3_io_hostInterface_cycle),
    .io_en(lsus_3_io_en),
    .io_in_0(lsus_3_io_in_0),
    .io_in_1(lsus_3_io_in_1),
    .io_out_0(lsus_3_io_out_0)
  );
  LSU_4 lsus_4 ( // @[CGRA.scala 364:21]
    .clock(lsus_4_clock),
    .reset(lsus_4_reset),
    .io_cfg_en(lsus_4_io_cfg_en),
    .io_cfg_addr(lsus_4_io_cfg_addr),
    .io_cfg_data(lsus_4_io_cfg_data),
    .io_hostInterface_read_addr(lsus_4_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_4_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_4_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_4_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_4_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_4_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_4_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_4_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_4_io_hostInterface_cycle),
    .io_en(lsus_4_io_en),
    .io_in_0(lsus_4_io_in_0),
    .io_in_1(lsus_4_io_in_1),
    .io_out_0(lsus_4_io_out_0)
  );
  LSU_5 lsus_5 ( // @[CGRA.scala 364:21]
    .clock(lsus_5_clock),
    .reset(lsus_5_reset),
    .io_cfg_en(lsus_5_io_cfg_en),
    .io_cfg_addr(lsus_5_io_cfg_addr),
    .io_cfg_data(lsus_5_io_cfg_data),
    .io_hostInterface_read_addr(lsus_5_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_5_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_5_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_5_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_5_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_5_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_5_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_5_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_5_io_hostInterface_cycle),
    .io_en(lsus_5_io_en),
    .io_in_0(lsus_5_io_in_0),
    .io_in_1(lsus_5_io_in_1),
    .io_out_0(lsus_5_io_out_0)
  );
  LSU_6 lsus_6 ( // @[CGRA.scala 364:21]
    .clock(lsus_6_clock),
    .reset(lsus_6_reset),
    .io_cfg_en(lsus_6_io_cfg_en),
    .io_cfg_addr(lsus_6_io_cfg_addr),
    .io_cfg_data(lsus_6_io_cfg_data),
    .io_hostInterface_read_addr(lsus_6_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_6_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_6_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_6_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_6_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_6_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_6_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_6_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_6_io_hostInterface_cycle),
    .io_en(lsus_6_io_en),
    .io_in_0(lsus_6_io_in_0),
    .io_in_1(lsus_6_io_in_1),
    .io_out_0(lsus_6_io_out_0)
  );
  LSU_7 lsus_7 ( // @[CGRA.scala 364:21]
    .clock(lsus_7_clock),
    .reset(lsus_7_reset),
    .io_cfg_en(lsus_7_io_cfg_en),
    .io_cfg_addr(lsus_7_io_cfg_addr),
    .io_cfg_data(lsus_7_io_cfg_data),
    .io_hostInterface_read_addr(lsus_7_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_7_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_7_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_7_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_7_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_7_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_7_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_7_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_7_io_hostInterface_cycle),
    .io_en(lsus_7_io_en),
    .io_in_0(lsus_7_io_in_0),
    .io_in_1(lsus_7_io_in_1),
    .io_out_0(lsus_7_io_out_0)
  );
  LSU_8 lsus_8 ( // @[CGRA.scala 364:21]
    .clock(lsus_8_clock),
    .reset(lsus_8_reset),
    .io_cfg_en(lsus_8_io_cfg_en),
    .io_cfg_addr(lsus_8_io_cfg_addr),
    .io_cfg_data(lsus_8_io_cfg_data),
    .io_hostInterface_read_addr(lsus_8_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_8_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_8_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_8_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_8_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_8_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_8_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_8_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_8_io_hostInterface_cycle),
    .io_en(lsus_8_io_en),
    .io_in_0(lsus_8_io_in_0),
    .io_in_1(lsus_8_io_in_1),
    .io_out_0(lsus_8_io_out_0)
  );
  LSU_9 lsus_9 ( // @[CGRA.scala 364:21]
    .clock(lsus_9_clock),
    .reset(lsus_9_reset),
    .io_cfg_en(lsus_9_io_cfg_en),
    .io_cfg_addr(lsus_9_io_cfg_addr),
    .io_cfg_data(lsus_9_io_cfg_data),
    .io_hostInterface_read_addr(lsus_9_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_9_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_9_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_9_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_9_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_9_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_9_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_9_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_9_io_hostInterface_cycle),
    .io_en(lsus_9_io_en),
    .io_in_0(lsus_9_io_in_0),
    .io_in_1(lsus_9_io_in_1),
    .io_out_0(lsus_9_io_out_0)
  );
  LSU_10 lsus_10 ( // @[CGRA.scala 364:21]
    .clock(lsus_10_clock),
    .reset(lsus_10_reset),
    .io_cfg_en(lsus_10_io_cfg_en),
    .io_cfg_addr(lsus_10_io_cfg_addr),
    .io_cfg_data(lsus_10_io_cfg_data),
    .io_hostInterface_read_addr(lsus_10_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_10_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_10_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_10_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_10_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_10_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_10_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_10_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_10_io_hostInterface_cycle),
    .io_en(lsus_10_io_en),
    .io_in_0(lsus_10_io_in_0),
    .io_in_1(lsus_10_io_in_1),
    .io_out_0(lsus_10_io_out_0)
  );
  LSU_11 lsus_11 ( // @[CGRA.scala 364:21]
    .clock(lsus_11_clock),
    .reset(lsus_11_reset),
    .io_cfg_en(lsus_11_io_cfg_en),
    .io_cfg_addr(lsus_11_io_cfg_addr),
    .io_cfg_data(lsus_11_io_cfg_data),
    .io_hostInterface_read_addr(lsus_11_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_11_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_11_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_11_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_11_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_11_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_11_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_11_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_11_io_hostInterface_cycle),
    .io_en(lsus_11_io_en),
    .io_in_0(lsus_11_io_in_0),
    .io_in_1(lsus_11_io_in_1),
    .io_out_0(lsus_11_io_out_0)
  );
  LSU_12 lsus_12 ( // @[CGRA.scala 364:21]
    .clock(lsus_12_clock),
    .reset(lsus_12_reset),
    .io_cfg_en(lsus_12_io_cfg_en),
    .io_cfg_addr(lsus_12_io_cfg_addr),
    .io_cfg_data(lsus_12_io_cfg_data),
    .io_hostInterface_read_addr(lsus_12_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_12_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_12_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_12_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_12_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_12_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_12_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_12_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_12_io_hostInterface_cycle),
    .io_en(lsus_12_io_en),
    .io_in_0(lsus_12_io_in_0),
    .io_in_1(lsus_12_io_in_1),
    .io_out_0(lsus_12_io_out_0)
  );
  LSU_13 lsus_13 ( // @[CGRA.scala 364:21]
    .clock(lsus_13_clock),
    .reset(lsus_13_reset),
    .io_cfg_en(lsus_13_io_cfg_en),
    .io_cfg_addr(lsus_13_io_cfg_addr),
    .io_cfg_data(lsus_13_io_cfg_data),
    .io_hostInterface_read_addr(lsus_13_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_13_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_13_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_13_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_13_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_13_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_13_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_13_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_13_io_hostInterface_cycle),
    .io_en(lsus_13_io_en),
    .io_in_0(lsus_13_io_in_0),
    .io_in_1(lsus_13_io_in_1),
    .io_out_0(lsus_13_io_out_0)
  );
  LSU_14 lsus_14 ( // @[CGRA.scala 364:21]
    .clock(lsus_14_clock),
    .reset(lsus_14_reset),
    .io_cfg_en(lsus_14_io_cfg_en),
    .io_cfg_addr(lsus_14_io_cfg_addr),
    .io_cfg_data(lsus_14_io_cfg_data),
    .io_hostInterface_read_addr(lsus_14_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_14_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_14_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_14_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_14_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_14_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_14_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_14_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_14_io_hostInterface_cycle),
    .io_en(lsus_14_io_en),
    .io_in_0(lsus_14_io_in_0),
    .io_in_1(lsus_14_io_in_1),
    .io_out_0(lsus_14_io_out_0)
  );
  LSU_15 lsus_15 ( // @[CGRA.scala 364:21]
    .clock(lsus_15_clock),
    .reset(lsus_15_reset),
    .io_cfg_en(lsus_15_io_cfg_en),
    .io_cfg_addr(lsus_15_io_cfg_addr),
    .io_cfg_data(lsus_15_io_cfg_data),
    .io_hostInterface_read_addr(lsus_15_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_15_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_15_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_15_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_15_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_15_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_15_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_15_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_15_io_hostInterface_cycle),
    .io_en(lsus_15_io_en),
    .io_in_0(lsus_15_io_in_0),
    .io_in_1(lsus_15_io_in_1),
    .io_out_0(lsus_15_io_out_0)
  );
  LSU_16 lsus_16 ( // @[CGRA.scala 364:21]
    .clock(lsus_16_clock),
    .reset(lsus_16_reset),
    .io_cfg_en(lsus_16_io_cfg_en),
    .io_cfg_addr(lsus_16_io_cfg_addr),
    .io_cfg_data(lsus_16_io_cfg_data),
    .io_hostInterface_read_addr(lsus_16_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_16_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_16_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_16_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_16_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_16_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_16_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_16_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_16_io_hostInterface_cycle),
    .io_en(lsus_16_io_en),
    .io_in_0(lsus_16_io_in_0),
    .io_in_1(lsus_16_io_in_1),
    .io_out_0(lsus_16_io_out_0)
  );
  LSU_17 lsus_17 ( // @[CGRA.scala 364:21]
    .clock(lsus_17_clock),
    .reset(lsus_17_reset),
    .io_cfg_en(lsus_17_io_cfg_en),
    .io_cfg_addr(lsus_17_io_cfg_addr),
    .io_cfg_data(lsus_17_io_cfg_data),
    .io_hostInterface_read_addr(lsus_17_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_17_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_17_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_17_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_17_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_17_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_17_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_17_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_17_io_hostInterface_cycle),
    .io_en(lsus_17_io_en),
    .io_in_0(lsus_17_io_in_0),
    .io_in_1(lsus_17_io_in_1),
    .io_out_0(lsus_17_io_out_0)
  );
  LSU_18 lsus_18 ( // @[CGRA.scala 364:21]
    .clock(lsus_18_clock),
    .reset(lsus_18_reset),
    .io_cfg_en(lsus_18_io_cfg_en),
    .io_cfg_addr(lsus_18_io_cfg_addr),
    .io_cfg_data(lsus_18_io_cfg_data),
    .io_hostInterface_read_addr(lsus_18_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_18_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_18_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_18_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_18_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_18_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_18_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_18_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_18_io_hostInterface_cycle),
    .io_en(lsus_18_io_en),
    .io_in_0(lsus_18_io_in_0),
    .io_in_1(lsus_18_io_in_1),
    .io_out_0(lsus_18_io_out_0)
  );
  LSU_19 lsus_19 ( // @[CGRA.scala 364:21]
    .clock(lsus_19_clock),
    .reset(lsus_19_reset),
    .io_cfg_en(lsus_19_io_cfg_en),
    .io_cfg_addr(lsus_19_io_cfg_addr),
    .io_cfg_data(lsus_19_io_cfg_data),
    .io_hostInterface_read_addr(lsus_19_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_19_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_19_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_19_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_19_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_19_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_19_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_19_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_19_io_hostInterface_cycle),
    .io_en(lsus_19_io_en),
    .io_in_0(lsus_19_io_in_0),
    .io_in_1(lsus_19_io_in_1),
    .io_out_0(lsus_19_io_out_0)
  );
  LSU_20 lsus_20 ( // @[CGRA.scala 364:21]
    .clock(lsus_20_clock),
    .reset(lsus_20_reset),
    .io_cfg_en(lsus_20_io_cfg_en),
    .io_cfg_addr(lsus_20_io_cfg_addr),
    .io_cfg_data(lsus_20_io_cfg_data),
    .io_hostInterface_read_addr(lsus_20_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_20_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_20_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_20_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_20_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_20_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_20_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_20_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_20_io_hostInterface_cycle),
    .io_en(lsus_20_io_en),
    .io_in_0(lsus_20_io_in_0),
    .io_in_1(lsus_20_io_in_1),
    .io_out_0(lsus_20_io_out_0)
  );
  LSU_21 lsus_21 ( // @[CGRA.scala 364:21]
    .clock(lsus_21_clock),
    .reset(lsus_21_reset),
    .io_cfg_en(lsus_21_io_cfg_en),
    .io_cfg_addr(lsus_21_io_cfg_addr),
    .io_cfg_data(lsus_21_io_cfg_data),
    .io_hostInterface_read_addr(lsus_21_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_21_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_21_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_21_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_21_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_21_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_21_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_21_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_21_io_hostInterface_cycle),
    .io_en(lsus_21_io_en),
    .io_in_0(lsus_21_io_in_0),
    .io_in_1(lsus_21_io_in_1),
    .io_out_0(lsus_21_io_out_0)
  );
  LSU_22 lsus_22 ( // @[CGRA.scala 364:21]
    .clock(lsus_22_clock),
    .reset(lsus_22_reset),
    .io_cfg_en(lsus_22_io_cfg_en),
    .io_cfg_addr(lsus_22_io_cfg_addr),
    .io_cfg_data(lsus_22_io_cfg_data),
    .io_hostInterface_read_addr(lsus_22_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_22_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_22_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_22_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_22_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_22_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_22_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_22_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_22_io_hostInterface_cycle),
    .io_en(lsus_22_io_en),
    .io_in_0(lsus_22_io_in_0),
    .io_in_1(lsus_22_io_in_1),
    .io_out_0(lsus_22_io_out_0)
  );
  LSU_23 lsus_23 ( // @[CGRA.scala 364:21]
    .clock(lsus_23_clock),
    .reset(lsus_23_reset),
    .io_cfg_en(lsus_23_io_cfg_en),
    .io_cfg_addr(lsus_23_io_cfg_addr),
    .io_cfg_data(lsus_23_io_cfg_data),
    .io_hostInterface_read_addr(lsus_23_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_23_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_23_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_23_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_23_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_23_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_23_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_23_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_23_io_hostInterface_cycle),
    .io_en(lsus_23_io_en),
    .io_in_0(lsus_23_io_in_0),
    .io_in_1(lsus_23_io_in_1),
    .io_out_0(lsus_23_io_out_0)
  );
  LSU_24 lsus_24 ( // @[CGRA.scala 364:21]
    .clock(lsus_24_clock),
    .reset(lsus_24_reset),
    .io_cfg_en(lsus_24_io_cfg_en),
    .io_cfg_addr(lsus_24_io_cfg_addr),
    .io_cfg_data(lsus_24_io_cfg_data),
    .io_hostInterface_read_addr(lsus_24_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_24_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_24_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_24_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_24_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_24_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_24_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_24_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_24_io_hostInterface_cycle),
    .io_en(lsus_24_io_en),
    .io_in_0(lsus_24_io_in_0),
    .io_in_1(lsus_24_io_in_1),
    .io_out_0(lsus_24_io_out_0)
  );
  LSU_25 lsus_25 ( // @[CGRA.scala 364:21]
    .clock(lsus_25_clock),
    .reset(lsus_25_reset),
    .io_cfg_en(lsus_25_io_cfg_en),
    .io_cfg_addr(lsus_25_io_cfg_addr),
    .io_cfg_data(lsus_25_io_cfg_data),
    .io_hostInterface_read_addr(lsus_25_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_25_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_25_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_25_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_25_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_25_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_25_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_25_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_25_io_hostInterface_cycle),
    .io_en(lsus_25_io_en),
    .io_in_0(lsus_25_io_in_0),
    .io_in_1(lsus_25_io_in_1),
    .io_out_0(lsus_25_io_out_0)
  );
  LSU_26 lsus_26 ( // @[CGRA.scala 364:21]
    .clock(lsus_26_clock),
    .reset(lsus_26_reset),
    .io_cfg_en(lsus_26_io_cfg_en),
    .io_cfg_addr(lsus_26_io_cfg_addr),
    .io_cfg_data(lsus_26_io_cfg_data),
    .io_hostInterface_read_addr(lsus_26_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_26_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_26_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_26_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_26_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_26_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_26_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_26_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_26_io_hostInterface_cycle),
    .io_en(lsus_26_io_en),
    .io_in_0(lsus_26_io_in_0),
    .io_in_1(lsus_26_io_in_1),
    .io_out_0(lsus_26_io_out_0)
  );
  LSU_27 lsus_27 ( // @[CGRA.scala 364:21]
    .clock(lsus_27_clock),
    .reset(lsus_27_reset),
    .io_cfg_en(lsus_27_io_cfg_en),
    .io_cfg_addr(lsus_27_io_cfg_addr),
    .io_cfg_data(lsus_27_io_cfg_data),
    .io_hostInterface_read_addr(lsus_27_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_27_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_27_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_27_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_27_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_27_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_27_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_27_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_27_io_hostInterface_cycle),
    .io_en(lsus_27_io_en),
    .io_in_0(lsus_27_io_in_0),
    .io_in_1(lsus_27_io_in_1),
    .io_out_0(lsus_27_io_out_0)
  );
  LSU_28 lsus_28 ( // @[CGRA.scala 364:21]
    .clock(lsus_28_clock),
    .reset(lsus_28_reset),
    .io_cfg_en(lsus_28_io_cfg_en),
    .io_cfg_addr(lsus_28_io_cfg_addr),
    .io_cfg_data(lsus_28_io_cfg_data),
    .io_hostInterface_read_addr(lsus_28_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_28_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_28_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_28_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_28_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_28_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_28_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_28_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_28_io_hostInterface_cycle),
    .io_en(lsus_28_io_en),
    .io_in_0(lsus_28_io_in_0),
    .io_in_1(lsus_28_io_in_1),
    .io_out_0(lsus_28_io_out_0)
  );
  LSU_29 lsus_29 ( // @[CGRA.scala 364:21]
    .clock(lsus_29_clock),
    .reset(lsus_29_reset),
    .io_cfg_en(lsus_29_io_cfg_en),
    .io_cfg_addr(lsus_29_io_cfg_addr),
    .io_cfg_data(lsus_29_io_cfg_data),
    .io_hostInterface_read_addr(lsus_29_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_29_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_29_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_29_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_29_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_29_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_29_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_29_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_29_io_hostInterface_cycle),
    .io_en(lsus_29_io_en),
    .io_in_0(lsus_29_io_in_0),
    .io_in_1(lsus_29_io_in_1),
    .io_out_0(lsus_29_io_out_0)
  );
  LSU_30 lsus_30 ( // @[CGRA.scala 364:21]
    .clock(lsus_30_clock),
    .reset(lsus_30_reset),
    .io_cfg_en(lsus_30_io_cfg_en),
    .io_cfg_addr(lsus_30_io_cfg_addr),
    .io_cfg_data(lsus_30_io_cfg_data),
    .io_hostInterface_read_addr(lsus_30_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_30_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_30_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_30_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_30_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_30_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_30_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_30_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_30_io_hostInterface_cycle),
    .io_en(lsus_30_io_en),
    .io_in_0(lsus_30_io_in_0),
    .io_in_1(lsus_30_io_in_1),
    .io_out_0(lsus_30_io_out_0)
  );
  LSU_31 lsus_31 ( // @[CGRA.scala 364:21]
    .clock(lsus_31_clock),
    .reset(lsus_31_reset),
    .io_cfg_en(lsus_31_io_cfg_en),
    .io_cfg_addr(lsus_31_io_cfg_addr),
    .io_cfg_data(lsus_31_io_cfg_data),
    .io_hostInterface_read_addr(lsus_31_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_31_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_31_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_31_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_31_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_31_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_31_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_31_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_31_io_hostInterface_cycle),
    .io_en(lsus_31_io_en),
    .io_in_0(lsus_31_io_in_0),
    .io_in_1(lsus_31_io_in_1),
    .io_out_0(lsus_31_io_out_0)
  );
  LSU_32 lsus_32 ( // @[CGRA.scala 364:21]
    .clock(lsus_32_clock),
    .reset(lsus_32_reset),
    .io_cfg_en(lsus_32_io_cfg_en),
    .io_cfg_addr(lsus_32_io_cfg_addr),
    .io_cfg_data(lsus_32_io_cfg_data),
    .io_hostInterface_read_addr(lsus_32_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_32_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_32_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_32_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_32_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_32_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_32_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_32_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_32_io_hostInterface_cycle),
    .io_en(lsus_32_io_en),
    .io_in_0(lsus_32_io_in_0),
    .io_in_1(lsus_32_io_in_1),
    .io_out_0(lsus_32_io_out_0)
  );
  LSU_33 lsus_33 ( // @[CGRA.scala 364:21]
    .clock(lsus_33_clock),
    .reset(lsus_33_reset),
    .io_cfg_en(lsus_33_io_cfg_en),
    .io_cfg_addr(lsus_33_io_cfg_addr),
    .io_cfg_data(lsus_33_io_cfg_data),
    .io_hostInterface_read_addr(lsus_33_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_33_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_33_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_33_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_33_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_33_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_33_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_33_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_33_io_hostInterface_cycle),
    .io_en(lsus_33_io_en),
    .io_in_0(lsus_33_io_in_0),
    .io_in_1(lsus_33_io_in_1),
    .io_out_0(lsus_33_io_out_0)
  );
  LSU_34 lsus_34 ( // @[CGRA.scala 364:21]
    .clock(lsus_34_clock),
    .reset(lsus_34_reset),
    .io_cfg_en(lsus_34_io_cfg_en),
    .io_cfg_addr(lsus_34_io_cfg_addr),
    .io_cfg_data(lsus_34_io_cfg_data),
    .io_hostInterface_read_addr(lsus_34_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_34_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_34_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_34_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_34_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_34_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_34_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_34_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_34_io_hostInterface_cycle),
    .io_en(lsus_34_io_en),
    .io_in_0(lsus_34_io_in_0),
    .io_in_1(lsus_34_io_in_1),
    .io_out_0(lsus_34_io_out_0)
  );
  LSU_35 lsus_35 ( // @[CGRA.scala 364:21]
    .clock(lsus_35_clock),
    .reset(lsus_35_reset),
    .io_cfg_en(lsus_35_io_cfg_en),
    .io_cfg_addr(lsus_35_io_cfg_addr),
    .io_cfg_data(lsus_35_io_cfg_data),
    .io_hostInterface_read_addr(lsus_35_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_35_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_35_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_35_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_35_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_35_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_35_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_35_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_35_io_hostInterface_cycle),
    .io_en(lsus_35_io_en),
    .io_in_0(lsus_35_io_in_0),
    .io_in_1(lsus_35_io_in_1),
    .io_out_0(lsus_35_io_out_0)
  );
  LSU_36 lsus_36 ( // @[CGRA.scala 364:21]
    .clock(lsus_36_clock),
    .reset(lsus_36_reset),
    .io_cfg_en(lsus_36_io_cfg_en),
    .io_cfg_addr(lsus_36_io_cfg_addr),
    .io_cfg_data(lsus_36_io_cfg_data),
    .io_hostInterface_read_addr(lsus_36_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_36_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_36_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_36_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_36_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_36_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_36_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_36_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_36_io_hostInterface_cycle),
    .io_en(lsus_36_io_en),
    .io_in_0(lsus_36_io_in_0),
    .io_in_1(lsus_36_io_in_1),
    .io_out_0(lsus_36_io_out_0)
  );
  LSU_37 lsus_37 ( // @[CGRA.scala 364:21]
    .clock(lsus_37_clock),
    .reset(lsus_37_reset),
    .io_cfg_en(lsus_37_io_cfg_en),
    .io_cfg_addr(lsus_37_io_cfg_addr),
    .io_cfg_data(lsus_37_io_cfg_data),
    .io_hostInterface_read_addr(lsus_37_io_hostInterface_read_addr),
    .io_hostInterface_read_data_ready(lsus_37_io_hostInterface_read_data_ready),
    .io_hostInterface_read_data_valid(lsus_37_io_hostInterface_read_data_valid),
    .io_hostInterface_read_data_bits(lsus_37_io_hostInterface_read_data_bits),
    .io_hostInterface_write_addr(lsus_37_io_hostInterface_write_addr),
    .io_hostInterface_write_data_ready(lsus_37_io_hostInterface_write_data_ready),
    .io_hostInterface_write_data_valid(lsus_37_io_hostInterface_write_data_valid),
    .io_hostInterface_write_data_bits(lsus_37_io_hostInterface_write_data_bits),
    .io_hostInterface_cycle(lsus_37_io_hostInterface_cycle),
    .io_en(lsus_37_io_en),
    .io_in_0(lsus_37_io_in_0),
    .io_in_1(lsus_37_io_in_1),
    .io_out_0(lsus_37_io_out_0)
  );
  assign io_hostInterface_0_read_data_valid = lsus_0_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_0_read_data_bits = lsus_0_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_0_write_data_ready = lsus_0_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_1_read_data_valid = lsus_1_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_1_read_data_bits = lsus_1_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_1_write_data_ready = lsus_1_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_2_read_data_valid = lsus_2_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_2_read_data_bits = lsus_2_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_2_write_data_ready = lsus_2_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_3_read_data_valid = lsus_3_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_3_read_data_bits = lsus_3_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_3_write_data_ready = lsus_3_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_4_read_data_valid = lsus_4_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_4_read_data_bits = lsus_4_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_4_write_data_ready = lsus_4_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_5_read_data_valid = lsus_5_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_5_read_data_bits = lsus_5_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_5_write_data_ready = lsus_5_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_6_read_data_valid = lsus_6_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_6_read_data_bits = lsus_6_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_6_write_data_ready = lsus_6_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_7_read_data_valid = lsus_7_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_7_read_data_bits = lsus_7_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_7_write_data_ready = lsus_7_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_8_read_data_valid = lsus_8_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_8_read_data_bits = lsus_8_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_8_write_data_ready = lsus_8_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_9_read_data_valid = lsus_9_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_9_read_data_bits = lsus_9_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_9_write_data_ready = lsus_9_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_10_read_data_valid = lsus_10_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_10_read_data_bits = lsus_10_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_10_write_data_ready = lsus_10_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_11_read_data_valid = lsus_11_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_11_read_data_bits = lsus_11_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_11_write_data_ready = lsus_11_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_12_read_data_valid = lsus_12_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_12_read_data_bits = lsus_12_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_12_write_data_ready = lsus_12_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_13_read_data_valid = lsus_13_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_13_read_data_bits = lsus_13_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_13_write_data_ready = lsus_13_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_14_read_data_valid = lsus_14_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_14_read_data_bits = lsus_14_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_14_write_data_ready = lsus_14_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_15_read_data_valid = lsus_15_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_15_read_data_bits = lsus_15_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_15_write_data_ready = lsus_15_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_16_read_data_valid = lsus_16_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_16_read_data_bits = lsus_16_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_16_write_data_ready = lsus_16_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_17_read_data_valid = lsus_17_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_17_read_data_bits = lsus_17_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_17_write_data_ready = lsus_17_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_18_read_data_valid = lsus_18_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_18_read_data_bits = lsus_18_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_18_write_data_ready = lsus_18_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_19_read_data_valid = lsus_19_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_19_read_data_bits = lsus_19_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_19_write_data_ready = lsus_19_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_20_read_data_valid = lsus_20_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_20_read_data_bits = lsus_20_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_20_write_data_ready = lsus_20_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_21_read_data_valid = lsus_21_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_21_read_data_bits = lsus_21_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_21_write_data_ready = lsus_21_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_22_read_data_valid = lsus_22_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_22_read_data_bits = lsus_22_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_22_write_data_ready = lsus_22_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_23_read_data_valid = lsus_23_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_23_read_data_bits = lsus_23_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_23_write_data_ready = lsus_23_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_24_read_data_valid = lsus_24_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_24_read_data_bits = lsus_24_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_24_write_data_ready = lsus_24_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_25_read_data_valid = lsus_25_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_25_read_data_bits = lsus_25_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_25_write_data_ready = lsus_25_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_26_read_data_valid = lsus_26_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_26_read_data_bits = lsus_26_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_26_write_data_ready = lsus_26_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_27_read_data_valid = lsus_27_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_27_read_data_bits = lsus_27_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_27_write_data_ready = lsus_27_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_28_read_data_valid = lsus_28_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_28_read_data_bits = lsus_28_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_28_write_data_ready = lsus_28_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_29_read_data_valid = lsus_29_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_29_read_data_bits = lsus_29_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_29_write_data_ready = lsus_29_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_30_read_data_valid = lsus_30_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_30_read_data_bits = lsus_30_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_30_write_data_ready = lsus_30_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_31_read_data_valid = lsus_31_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_31_read_data_bits = lsus_31_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_31_write_data_ready = lsus_31_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_32_read_data_valid = lsus_32_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_32_read_data_bits = lsus_32_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_32_write_data_ready = lsus_32_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_33_read_data_valid = lsus_33_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_33_read_data_bits = lsus_33_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_33_write_data_ready = lsus_33_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_34_read_data_valid = lsus_34_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_34_read_data_bits = lsus_34_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_34_write_data_ready = lsus_34_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_35_read_data_valid = lsus_35_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_35_read_data_bits = lsus_35_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_35_write_data_ready = lsus_35_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_36_read_data_valid = lsus_36_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_36_read_data_bits = lsus_36_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_36_write_data_ready = lsus_36_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_hostInterface_37_read_data_valid = lsus_37_io_hostInterface_read_data_valid; // @[CGRA.scala 595:36]
  assign io_hostInterface_37_read_data_bits = lsus_37_io_hostInterface_read_data_bits; // @[CGRA.scala 595:36]
  assign io_hostInterface_37_write_data_ready = lsus_37_io_hostInterface_write_data_ready; // @[CGRA.scala 595:36]
  assign io_out_0 = obs_0_io_out_0; // @[CGRA.scala 443:26]
  assign io_out_1 = obs_1_io_out_0; // @[CGRA.scala 443:26]
  assign io_out_2 = obs_2_io_out_0; // @[CGRA.scala 443:26]
  assign io_out_3 = obs_3_io_out_0; // @[CGRA.scala 443:26]
  assign io_out_4 = obs_4_io_out_0; // @[CGRA.scala 443:26]
  assign io_out_5 = obs_5_io_out_0; // @[CGRA.scala 443:26]
  assign ibs_0_io_in_0 = io_in_0; // @[CGRA.scala 414:19]
  assign ibs_1_io_in_0 = io_in_1; // @[CGRA.scala 414:19]
  assign ibs_2_io_in_0 = io_in_2; // @[CGRA.scala 414:19]
  assign ibs_3_io_in_0 = io_in_3; // @[CGRA.scala 414:19]
  assign ibs_4_io_in_0 = io_in_4; // @[CGRA.scala 414:19]
  assign ibs_5_io_in_0 = io_in_5; // @[CGRA.scala 414:19]
  assign obs_0_clock = clock;
  assign obs_0_reset = reset;
  assign obs_0_io_cfg_en = cfgRegs_0[46]; // @[CGRA.scala 652:24]
  assign obs_0_io_cfg_addr = cfgRegs_0[45:32]; // @[CGRA.scala 653:24]
  assign obs_0_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 654:24]
  assign obs_0_io_in_0 = gibs_0_io_ipinNE_0; // @[CGRA.scala 450:14]
  assign obs_0_io_in_1 = gibs_1_io_ipinNW_0; // @[CGRA.scala 454:14]
  assign obs_1_clock = clock;
  assign obs_1_reset = reset;
  assign obs_1_io_cfg_en = cfgRegs_0[46]; // @[CGRA.scala 652:24]
  assign obs_1_io_cfg_addr = cfgRegs_0[45:32]; // @[CGRA.scala 653:24]
  assign obs_1_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 654:24]
  assign obs_1_io_in_0 = gibs_1_io_ipinNE_0; // @[CGRA.scala 450:14]
  assign obs_1_io_in_1 = gibs_2_io_ipinNW_0; // @[CGRA.scala 454:14]
  assign obs_2_clock = clock;
  assign obs_2_reset = reset;
  assign obs_2_io_cfg_en = cfgRegs_0[46]; // @[CGRA.scala 652:24]
  assign obs_2_io_cfg_addr = cfgRegs_0[45:32]; // @[CGRA.scala 653:24]
  assign obs_2_io_cfg_data = cfgRegs_0[31:0]; // @[CGRA.scala 654:24]
  assign obs_2_io_in_0 = gibs_2_io_ipinNE_0; // @[CGRA.scala 450:14]
  assign obs_2_io_in_1 = gibs_3_io_ipinNW_0; // @[CGRA.scala 454:14]
  assign obs_3_clock = clock;
  assign obs_3_reset = reset;
  assign obs_3_io_cfg_en = cfgRegs_41[46]; // @[CGRA.scala 661:26]
  assign obs_3_io_cfg_addr = cfgRegs_41[45:32]; // @[CGRA.scala 662:26]
  assign obs_3_io_cfg_data = cfgRegs_41[31:0]; // @[CGRA.scala 663:26]
  assign obs_3_io_in_0 = gibs_76_io_ipinSE_0; // @[CGRA.scala 461:14]
  assign obs_3_io_in_1 = gibs_77_io_ipinSW_0; // @[CGRA.scala 465:14]
  assign obs_4_clock = clock;
  assign obs_4_reset = reset;
  assign obs_4_io_cfg_en = cfgRegs_41[46]; // @[CGRA.scala 661:26]
  assign obs_4_io_cfg_addr = cfgRegs_41[45:32]; // @[CGRA.scala 662:26]
  assign obs_4_io_cfg_data = cfgRegs_41[31:0]; // @[CGRA.scala 663:26]
  assign obs_4_io_in_0 = gibs_77_io_ipinSE_0; // @[CGRA.scala 461:14]
  assign obs_4_io_in_1 = gibs_78_io_ipinSW_0; // @[CGRA.scala 465:14]
  assign obs_5_clock = clock;
  assign obs_5_reset = reset;
  assign obs_5_io_cfg_en = cfgRegs_41[46]; // @[CGRA.scala 661:26]
  assign obs_5_io_cfg_addr = cfgRegs_41[45:32]; // @[CGRA.scala 662:26]
  assign obs_5_io_cfg_data = cfgRegs_41[31:0]; // @[CGRA.scala 663:26]
  assign obs_5_io_in_0 = gibs_78_io_ipinSE_0; // @[CGRA.scala 461:14]
  assign obs_5_io_in_1 = gibs_79_io_ipinSW_0; // @[CGRA.scala 465:14]
  assign pes_0_clock = clock;
  assign pes_0_reset = reset;
  assign pes_0_io_cfg_en = cfgRegs_2[46]; // @[CGRA.scala 671:37]
  assign pes_0_io_cfg_addr = cfgRegs_2[45:32]; // @[CGRA.scala 672:39]
  assign pes_0_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 673:39]
  assign pes_0_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_0_io_in_0 = gibs_0_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_0_io_in_1 = gibs_1_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_0_io_in_2 = gibs_4_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_0_io_in_3 = gibs_5_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_0_io_in_4 = gibs_0_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_0_io_in_5 = gibs_1_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_0_io_in_6 = gibs_4_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_0_io_in_7 = gibs_5_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_1_clock = clock;
  assign pes_1_reset = reset;
  assign pes_1_io_cfg_en = cfgRegs_2[46]; // @[CGRA.scala 671:37]
  assign pes_1_io_cfg_addr = cfgRegs_2[45:32]; // @[CGRA.scala 672:39]
  assign pes_1_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 673:39]
  assign pes_1_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_1_io_in_0 = gibs_1_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_1_io_in_1 = gibs_2_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_1_io_in_2 = gibs_5_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_1_io_in_3 = gibs_6_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_1_io_in_4 = gibs_1_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_1_io_in_5 = gibs_2_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_1_io_in_6 = gibs_5_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_1_io_in_7 = gibs_6_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_2_clock = clock;
  assign pes_2_reset = reset;
  assign pes_2_io_cfg_en = cfgRegs_2[46]; // @[CGRA.scala 671:37]
  assign pes_2_io_cfg_addr = cfgRegs_2[45:32]; // @[CGRA.scala 672:39]
  assign pes_2_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 673:39]
  assign pes_2_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_2_io_in_0 = gibs_2_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_2_io_in_1 = gibs_3_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_2_io_in_2 = gibs_6_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_2_io_in_3 = gibs_7_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_2_io_in_4 = gibs_2_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_2_io_in_5 = gibs_3_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_2_io_in_6 = gibs_6_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_2_io_in_7 = gibs_7_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_3_clock = clock;
  assign pes_3_reset = reset;
  assign pes_3_io_cfg_en = cfgRegs_4[46]; // @[CGRA.scala 671:37]
  assign pes_3_io_cfg_addr = cfgRegs_4[45:32]; // @[CGRA.scala 672:39]
  assign pes_3_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 673:39]
  assign pes_3_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_3_io_in_0 = gibs_4_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_3_io_in_1 = gibs_5_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_3_io_in_2 = gibs_8_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_3_io_in_3 = gibs_9_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_3_io_in_4 = gibs_4_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_3_io_in_5 = gibs_5_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_3_io_in_6 = gibs_8_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_3_io_in_7 = gibs_9_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_4_clock = clock;
  assign pes_4_reset = reset;
  assign pes_4_io_cfg_en = cfgRegs_4[46]; // @[CGRA.scala 671:37]
  assign pes_4_io_cfg_addr = cfgRegs_4[45:32]; // @[CGRA.scala 672:39]
  assign pes_4_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 673:39]
  assign pes_4_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_4_io_in_0 = gibs_5_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_4_io_in_1 = gibs_6_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_4_io_in_2 = gibs_9_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_4_io_in_3 = gibs_10_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_4_io_in_4 = gibs_5_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_4_io_in_5 = gibs_6_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_4_io_in_6 = gibs_9_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_4_io_in_7 = gibs_10_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_5_clock = clock;
  assign pes_5_reset = reset;
  assign pes_5_io_cfg_en = cfgRegs_4[46]; // @[CGRA.scala 671:37]
  assign pes_5_io_cfg_addr = cfgRegs_4[45:32]; // @[CGRA.scala 672:39]
  assign pes_5_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 673:39]
  assign pes_5_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_5_io_in_0 = gibs_6_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_5_io_in_1 = gibs_7_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_5_io_in_2 = gibs_10_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_5_io_in_3 = gibs_11_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_5_io_in_4 = gibs_6_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_5_io_in_5 = gibs_7_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_5_io_in_6 = gibs_10_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_5_io_in_7 = gibs_11_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_6_clock = clock;
  assign pes_6_reset = reset;
  assign pes_6_io_cfg_en = cfgRegs_6[46]; // @[CGRA.scala 671:37]
  assign pes_6_io_cfg_addr = cfgRegs_6[45:32]; // @[CGRA.scala 672:39]
  assign pes_6_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 673:39]
  assign pes_6_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_6_io_in_0 = gibs_8_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_6_io_in_1 = gibs_9_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_6_io_in_2 = gibs_12_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_6_io_in_3 = gibs_13_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_6_io_in_4 = gibs_8_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_6_io_in_5 = gibs_9_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_6_io_in_6 = gibs_12_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_6_io_in_7 = gibs_13_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_7_clock = clock;
  assign pes_7_reset = reset;
  assign pes_7_io_cfg_en = cfgRegs_6[46]; // @[CGRA.scala 671:37]
  assign pes_7_io_cfg_addr = cfgRegs_6[45:32]; // @[CGRA.scala 672:39]
  assign pes_7_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 673:39]
  assign pes_7_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_7_io_in_0 = gibs_9_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_7_io_in_1 = gibs_10_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_7_io_in_2 = gibs_13_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_7_io_in_3 = gibs_14_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_7_io_in_4 = gibs_9_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_7_io_in_5 = gibs_10_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_7_io_in_6 = gibs_13_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_7_io_in_7 = gibs_14_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_8_clock = clock;
  assign pes_8_reset = reset;
  assign pes_8_io_cfg_en = cfgRegs_6[46]; // @[CGRA.scala 671:37]
  assign pes_8_io_cfg_addr = cfgRegs_6[45:32]; // @[CGRA.scala 672:39]
  assign pes_8_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 673:39]
  assign pes_8_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_8_io_in_0 = gibs_10_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_8_io_in_1 = gibs_11_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_8_io_in_2 = gibs_14_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_8_io_in_3 = gibs_15_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_8_io_in_4 = gibs_10_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_8_io_in_5 = gibs_11_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_8_io_in_6 = gibs_14_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_8_io_in_7 = gibs_15_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_9_clock = clock;
  assign pes_9_reset = reset;
  assign pes_9_io_cfg_en = cfgRegs_8[46]; // @[CGRA.scala 671:37]
  assign pes_9_io_cfg_addr = cfgRegs_8[45:32]; // @[CGRA.scala 672:39]
  assign pes_9_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 673:39]
  assign pes_9_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_9_io_in_0 = gibs_12_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_9_io_in_1 = gibs_13_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_9_io_in_2 = gibs_16_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_9_io_in_3 = gibs_17_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_9_io_in_4 = gibs_12_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_9_io_in_5 = gibs_13_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_9_io_in_6 = gibs_16_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_9_io_in_7 = gibs_17_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_10_clock = clock;
  assign pes_10_reset = reset;
  assign pes_10_io_cfg_en = cfgRegs_8[46]; // @[CGRA.scala 671:37]
  assign pes_10_io_cfg_addr = cfgRegs_8[45:32]; // @[CGRA.scala 672:39]
  assign pes_10_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 673:39]
  assign pes_10_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_10_io_in_0 = gibs_13_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_10_io_in_1 = gibs_14_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_10_io_in_2 = gibs_17_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_10_io_in_3 = gibs_18_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_10_io_in_4 = gibs_13_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_10_io_in_5 = gibs_14_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_10_io_in_6 = gibs_17_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_10_io_in_7 = gibs_18_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_11_clock = clock;
  assign pes_11_reset = reset;
  assign pes_11_io_cfg_en = cfgRegs_8[46]; // @[CGRA.scala 671:37]
  assign pes_11_io_cfg_addr = cfgRegs_8[45:32]; // @[CGRA.scala 672:39]
  assign pes_11_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 673:39]
  assign pes_11_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_11_io_in_0 = gibs_14_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_11_io_in_1 = gibs_15_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_11_io_in_2 = gibs_18_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_11_io_in_3 = gibs_19_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_11_io_in_4 = gibs_14_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_11_io_in_5 = gibs_15_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_11_io_in_6 = gibs_18_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_11_io_in_7 = gibs_19_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_12_clock = clock;
  assign pes_12_reset = reset;
  assign pes_12_io_cfg_en = cfgRegs_10[46]; // @[CGRA.scala 671:37]
  assign pes_12_io_cfg_addr = cfgRegs_10[45:32]; // @[CGRA.scala 672:39]
  assign pes_12_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 673:39]
  assign pes_12_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_12_io_in_0 = gibs_16_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_12_io_in_1 = gibs_17_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_12_io_in_2 = gibs_20_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_12_io_in_3 = gibs_21_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_12_io_in_4 = gibs_16_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_12_io_in_5 = gibs_17_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_12_io_in_6 = gibs_20_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_12_io_in_7 = gibs_21_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_13_clock = clock;
  assign pes_13_reset = reset;
  assign pes_13_io_cfg_en = cfgRegs_10[46]; // @[CGRA.scala 671:37]
  assign pes_13_io_cfg_addr = cfgRegs_10[45:32]; // @[CGRA.scala 672:39]
  assign pes_13_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 673:39]
  assign pes_13_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_13_io_in_0 = gibs_17_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_13_io_in_1 = gibs_18_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_13_io_in_2 = gibs_21_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_13_io_in_3 = gibs_22_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_13_io_in_4 = gibs_17_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_13_io_in_5 = gibs_18_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_13_io_in_6 = gibs_21_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_13_io_in_7 = gibs_22_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_14_clock = clock;
  assign pes_14_reset = reset;
  assign pes_14_io_cfg_en = cfgRegs_10[46]; // @[CGRA.scala 671:37]
  assign pes_14_io_cfg_addr = cfgRegs_10[45:32]; // @[CGRA.scala 672:39]
  assign pes_14_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 673:39]
  assign pes_14_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_14_io_in_0 = gibs_18_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_14_io_in_1 = gibs_19_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_14_io_in_2 = gibs_22_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_14_io_in_3 = gibs_23_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_14_io_in_4 = gibs_18_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_14_io_in_5 = gibs_19_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_14_io_in_6 = gibs_22_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_14_io_in_7 = gibs_23_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_15_clock = clock;
  assign pes_15_reset = reset;
  assign pes_15_io_cfg_en = cfgRegs_12[46]; // @[CGRA.scala 671:37]
  assign pes_15_io_cfg_addr = cfgRegs_12[45:32]; // @[CGRA.scala 672:39]
  assign pes_15_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 673:39]
  assign pes_15_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_15_io_in_0 = gibs_20_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_15_io_in_1 = gibs_21_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_15_io_in_2 = gibs_24_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_15_io_in_3 = gibs_25_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_15_io_in_4 = gibs_20_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_15_io_in_5 = gibs_21_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_15_io_in_6 = gibs_24_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_15_io_in_7 = gibs_25_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_16_clock = clock;
  assign pes_16_reset = reset;
  assign pes_16_io_cfg_en = cfgRegs_12[46]; // @[CGRA.scala 671:37]
  assign pes_16_io_cfg_addr = cfgRegs_12[45:32]; // @[CGRA.scala 672:39]
  assign pes_16_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 673:39]
  assign pes_16_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_16_io_in_0 = gibs_21_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_16_io_in_1 = gibs_22_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_16_io_in_2 = gibs_25_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_16_io_in_3 = gibs_26_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_16_io_in_4 = gibs_21_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_16_io_in_5 = gibs_22_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_16_io_in_6 = gibs_25_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_16_io_in_7 = gibs_26_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_17_clock = clock;
  assign pes_17_reset = reset;
  assign pes_17_io_cfg_en = cfgRegs_12[46]; // @[CGRA.scala 671:37]
  assign pes_17_io_cfg_addr = cfgRegs_12[45:32]; // @[CGRA.scala 672:39]
  assign pes_17_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 673:39]
  assign pes_17_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_17_io_in_0 = gibs_22_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_17_io_in_1 = gibs_23_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_17_io_in_2 = gibs_26_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_17_io_in_3 = gibs_27_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_17_io_in_4 = gibs_22_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_17_io_in_5 = gibs_23_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_17_io_in_6 = gibs_26_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_17_io_in_7 = gibs_27_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_18_clock = clock;
  assign pes_18_reset = reset;
  assign pes_18_io_cfg_en = cfgRegs_14[46]; // @[CGRA.scala 671:37]
  assign pes_18_io_cfg_addr = cfgRegs_14[45:32]; // @[CGRA.scala 672:39]
  assign pes_18_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 673:39]
  assign pes_18_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_18_io_in_0 = gibs_24_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_18_io_in_1 = gibs_25_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_18_io_in_2 = gibs_28_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_18_io_in_3 = gibs_29_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_18_io_in_4 = gibs_24_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_18_io_in_5 = gibs_25_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_18_io_in_6 = gibs_28_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_18_io_in_7 = gibs_29_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_19_clock = clock;
  assign pes_19_reset = reset;
  assign pes_19_io_cfg_en = cfgRegs_14[46]; // @[CGRA.scala 671:37]
  assign pes_19_io_cfg_addr = cfgRegs_14[45:32]; // @[CGRA.scala 672:39]
  assign pes_19_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 673:39]
  assign pes_19_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_19_io_in_0 = gibs_25_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_19_io_in_1 = gibs_26_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_19_io_in_2 = gibs_29_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_19_io_in_3 = gibs_30_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_19_io_in_4 = gibs_25_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_19_io_in_5 = gibs_26_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_19_io_in_6 = gibs_29_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_19_io_in_7 = gibs_30_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_20_clock = clock;
  assign pes_20_reset = reset;
  assign pes_20_io_cfg_en = cfgRegs_14[46]; // @[CGRA.scala 671:37]
  assign pes_20_io_cfg_addr = cfgRegs_14[45:32]; // @[CGRA.scala 672:39]
  assign pes_20_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 673:39]
  assign pes_20_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_20_io_in_0 = gibs_26_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_20_io_in_1 = gibs_27_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_20_io_in_2 = gibs_30_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_20_io_in_3 = gibs_31_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_20_io_in_4 = gibs_26_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_20_io_in_5 = gibs_27_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_20_io_in_6 = gibs_30_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_20_io_in_7 = gibs_31_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_21_clock = clock;
  assign pes_21_reset = reset;
  assign pes_21_io_cfg_en = cfgRegs_16[46]; // @[CGRA.scala 671:37]
  assign pes_21_io_cfg_addr = cfgRegs_16[45:32]; // @[CGRA.scala 672:39]
  assign pes_21_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 673:39]
  assign pes_21_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_21_io_in_0 = gibs_28_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_21_io_in_1 = gibs_29_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_21_io_in_2 = gibs_32_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_21_io_in_3 = gibs_33_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_21_io_in_4 = gibs_28_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_21_io_in_5 = gibs_29_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_21_io_in_6 = gibs_32_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_21_io_in_7 = gibs_33_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_22_clock = clock;
  assign pes_22_reset = reset;
  assign pes_22_io_cfg_en = cfgRegs_16[46]; // @[CGRA.scala 671:37]
  assign pes_22_io_cfg_addr = cfgRegs_16[45:32]; // @[CGRA.scala 672:39]
  assign pes_22_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 673:39]
  assign pes_22_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_22_io_in_0 = gibs_29_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_22_io_in_1 = gibs_30_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_22_io_in_2 = gibs_33_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_22_io_in_3 = gibs_34_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_22_io_in_4 = gibs_29_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_22_io_in_5 = gibs_30_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_22_io_in_6 = gibs_33_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_22_io_in_7 = gibs_34_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_23_clock = clock;
  assign pes_23_reset = reset;
  assign pes_23_io_cfg_en = cfgRegs_16[46]; // @[CGRA.scala 671:37]
  assign pes_23_io_cfg_addr = cfgRegs_16[45:32]; // @[CGRA.scala 672:39]
  assign pes_23_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 673:39]
  assign pes_23_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_23_io_in_0 = gibs_30_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_23_io_in_1 = gibs_31_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_23_io_in_2 = gibs_34_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_23_io_in_3 = gibs_35_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_23_io_in_4 = gibs_30_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_23_io_in_5 = gibs_31_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_23_io_in_6 = gibs_34_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_23_io_in_7 = gibs_35_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_24_clock = clock;
  assign pes_24_reset = reset;
  assign pes_24_io_cfg_en = cfgRegs_18[46]; // @[CGRA.scala 671:37]
  assign pes_24_io_cfg_addr = cfgRegs_18[45:32]; // @[CGRA.scala 672:39]
  assign pes_24_io_cfg_data = cfgRegs_18[31:0]; // @[CGRA.scala 673:39]
  assign pes_24_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_24_io_in_0 = gibs_32_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_24_io_in_1 = gibs_33_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_24_io_in_2 = gibs_36_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_24_io_in_3 = gibs_37_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_24_io_in_4 = gibs_32_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_24_io_in_5 = gibs_33_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_24_io_in_6 = gibs_36_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_24_io_in_7 = gibs_37_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_25_clock = clock;
  assign pes_25_reset = reset;
  assign pes_25_io_cfg_en = cfgRegs_18[46]; // @[CGRA.scala 671:37]
  assign pes_25_io_cfg_addr = cfgRegs_18[45:32]; // @[CGRA.scala 672:39]
  assign pes_25_io_cfg_data = cfgRegs_18[31:0]; // @[CGRA.scala 673:39]
  assign pes_25_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_25_io_in_0 = gibs_33_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_25_io_in_1 = gibs_34_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_25_io_in_2 = gibs_37_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_25_io_in_3 = gibs_38_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_25_io_in_4 = gibs_33_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_25_io_in_5 = gibs_34_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_25_io_in_6 = gibs_37_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_25_io_in_7 = gibs_38_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_26_clock = clock;
  assign pes_26_reset = reset;
  assign pes_26_io_cfg_en = cfgRegs_18[46]; // @[CGRA.scala 671:37]
  assign pes_26_io_cfg_addr = cfgRegs_18[45:32]; // @[CGRA.scala 672:39]
  assign pes_26_io_cfg_data = cfgRegs_18[31:0]; // @[CGRA.scala 673:39]
  assign pes_26_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_26_io_in_0 = gibs_34_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_26_io_in_1 = gibs_35_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_26_io_in_2 = gibs_38_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_26_io_in_3 = gibs_39_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_26_io_in_4 = gibs_34_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_26_io_in_5 = gibs_35_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_26_io_in_6 = gibs_38_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_26_io_in_7 = gibs_39_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_27_clock = clock;
  assign pes_27_reset = reset;
  assign pes_27_io_cfg_en = cfgRegs_20[46]; // @[CGRA.scala 671:37]
  assign pes_27_io_cfg_addr = cfgRegs_20[45:32]; // @[CGRA.scala 672:39]
  assign pes_27_io_cfg_data = cfgRegs_20[31:0]; // @[CGRA.scala 673:39]
  assign pes_27_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_27_io_in_0 = gibs_36_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_27_io_in_1 = gibs_37_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_27_io_in_2 = gibs_40_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_27_io_in_3 = gibs_41_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_27_io_in_4 = gibs_36_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_27_io_in_5 = gibs_37_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_27_io_in_6 = gibs_40_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_27_io_in_7 = gibs_41_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_28_clock = clock;
  assign pes_28_reset = reset;
  assign pes_28_io_cfg_en = cfgRegs_20[46]; // @[CGRA.scala 671:37]
  assign pes_28_io_cfg_addr = cfgRegs_20[45:32]; // @[CGRA.scala 672:39]
  assign pes_28_io_cfg_data = cfgRegs_20[31:0]; // @[CGRA.scala 673:39]
  assign pes_28_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_28_io_in_0 = gibs_37_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_28_io_in_1 = gibs_38_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_28_io_in_2 = gibs_41_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_28_io_in_3 = gibs_42_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_28_io_in_4 = gibs_37_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_28_io_in_5 = gibs_38_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_28_io_in_6 = gibs_41_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_28_io_in_7 = gibs_42_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_29_clock = clock;
  assign pes_29_reset = reset;
  assign pes_29_io_cfg_en = cfgRegs_20[46]; // @[CGRA.scala 671:37]
  assign pes_29_io_cfg_addr = cfgRegs_20[45:32]; // @[CGRA.scala 672:39]
  assign pes_29_io_cfg_data = cfgRegs_20[31:0]; // @[CGRA.scala 673:39]
  assign pes_29_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_29_io_in_0 = gibs_38_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_29_io_in_1 = gibs_39_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_29_io_in_2 = gibs_42_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_29_io_in_3 = gibs_43_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_29_io_in_4 = gibs_38_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_29_io_in_5 = gibs_39_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_29_io_in_6 = gibs_42_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_29_io_in_7 = gibs_43_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_30_clock = clock;
  assign pes_30_reset = reset;
  assign pes_30_io_cfg_en = cfgRegs_22[46]; // @[CGRA.scala 671:37]
  assign pes_30_io_cfg_addr = cfgRegs_22[45:32]; // @[CGRA.scala 672:39]
  assign pes_30_io_cfg_data = cfgRegs_22[31:0]; // @[CGRA.scala 673:39]
  assign pes_30_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_30_io_in_0 = gibs_40_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_30_io_in_1 = gibs_41_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_30_io_in_2 = gibs_44_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_30_io_in_3 = gibs_45_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_30_io_in_4 = gibs_40_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_30_io_in_5 = gibs_41_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_30_io_in_6 = gibs_44_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_30_io_in_7 = gibs_45_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_31_clock = clock;
  assign pes_31_reset = reset;
  assign pes_31_io_cfg_en = cfgRegs_22[46]; // @[CGRA.scala 671:37]
  assign pes_31_io_cfg_addr = cfgRegs_22[45:32]; // @[CGRA.scala 672:39]
  assign pes_31_io_cfg_data = cfgRegs_22[31:0]; // @[CGRA.scala 673:39]
  assign pes_31_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_31_io_in_0 = gibs_41_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_31_io_in_1 = gibs_42_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_31_io_in_2 = gibs_45_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_31_io_in_3 = gibs_46_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_31_io_in_4 = gibs_41_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_31_io_in_5 = gibs_42_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_31_io_in_6 = gibs_45_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_31_io_in_7 = gibs_46_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_32_clock = clock;
  assign pes_32_reset = reset;
  assign pes_32_io_cfg_en = cfgRegs_22[46]; // @[CGRA.scala 671:37]
  assign pes_32_io_cfg_addr = cfgRegs_22[45:32]; // @[CGRA.scala 672:39]
  assign pes_32_io_cfg_data = cfgRegs_22[31:0]; // @[CGRA.scala 673:39]
  assign pes_32_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_32_io_in_0 = gibs_42_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_32_io_in_1 = gibs_43_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_32_io_in_2 = gibs_46_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_32_io_in_3 = gibs_47_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_32_io_in_4 = gibs_42_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_32_io_in_5 = gibs_43_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_32_io_in_6 = gibs_46_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_32_io_in_7 = gibs_47_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_33_clock = clock;
  assign pes_33_reset = reset;
  assign pes_33_io_cfg_en = cfgRegs_24[46]; // @[CGRA.scala 671:37]
  assign pes_33_io_cfg_addr = cfgRegs_24[45:32]; // @[CGRA.scala 672:39]
  assign pes_33_io_cfg_data = cfgRegs_24[31:0]; // @[CGRA.scala 673:39]
  assign pes_33_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_33_io_in_0 = gibs_44_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_33_io_in_1 = gibs_45_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_33_io_in_2 = gibs_48_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_33_io_in_3 = gibs_49_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_33_io_in_4 = gibs_44_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_33_io_in_5 = gibs_45_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_33_io_in_6 = gibs_48_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_33_io_in_7 = gibs_49_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_34_clock = clock;
  assign pes_34_reset = reset;
  assign pes_34_io_cfg_en = cfgRegs_24[46]; // @[CGRA.scala 671:37]
  assign pes_34_io_cfg_addr = cfgRegs_24[45:32]; // @[CGRA.scala 672:39]
  assign pes_34_io_cfg_data = cfgRegs_24[31:0]; // @[CGRA.scala 673:39]
  assign pes_34_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_34_io_in_0 = gibs_45_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_34_io_in_1 = gibs_46_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_34_io_in_2 = gibs_49_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_34_io_in_3 = gibs_50_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_34_io_in_4 = gibs_45_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_34_io_in_5 = gibs_46_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_34_io_in_6 = gibs_49_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_34_io_in_7 = gibs_50_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_35_clock = clock;
  assign pes_35_reset = reset;
  assign pes_35_io_cfg_en = cfgRegs_24[46]; // @[CGRA.scala 671:37]
  assign pes_35_io_cfg_addr = cfgRegs_24[45:32]; // @[CGRA.scala 672:39]
  assign pes_35_io_cfg_data = cfgRegs_24[31:0]; // @[CGRA.scala 673:39]
  assign pes_35_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_35_io_in_0 = gibs_46_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_35_io_in_1 = gibs_47_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_35_io_in_2 = gibs_50_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_35_io_in_3 = gibs_51_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_35_io_in_4 = gibs_46_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_35_io_in_5 = gibs_47_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_35_io_in_6 = gibs_50_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_35_io_in_7 = gibs_51_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_36_clock = clock;
  assign pes_36_reset = reset;
  assign pes_36_io_cfg_en = cfgRegs_26[46]; // @[CGRA.scala 671:37]
  assign pes_36_io_cfg_addr = cfgRegs_26[45:32]; // @[CGRA.scala 672:39]
  assign pes_36_io_cfg_data = cfgRegs_26[31:0]; // @[CGRA.scala 673:39]
  assign pes_36_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_36_io_in_0 = gibs_48_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_36_io_in_1 = gibs_49_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_36_io_in_2 = gibs_52_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_36_io_in_3 = gibs_53_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_36_io_in_4 = gibs_48_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_36_io_in_5 = gibs_49_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_36_io_in_6 = gibs_52_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_36_io_in_7 = gibs_53_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_37_clock = clock;
  assign pes_37_reset = reset;
  assign pes_37_io_cfg_en = cfgRegs_26[46]; // @[CGRA.scala 671:37]
  assign pes_37_io_cfg_addr = cfgRegs_26[45:32]; // @[CGRA.scala 672:39]
  assign pes_37_io_cfg_data = cfgRegs_26[31:0]; // @[CGRA.scala 673:39]
  assign pes_37_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_37_io_in_0 = gibs_49_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_37_io_in_1 = gibs_50_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_37_io_in_2 = gibs_53_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_37_io_in_3 = gibs_54_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_37_io_in_4 = gibs_49_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_37_io_in_5 = gibs_50_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_37_io_in_6 = gibs_53_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_37_io_in_7 = gibs_54_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_38_clock = clock;
  assign pes_38_reset = reset;
  assign pes_38_io_cfg_en = cfgRegs_26[46]; // @[CGRA.scala 671:37]
  assign pes_38_io_cfg_addr = cfgRegs_26[45:32]; // @[CGRA.scala 672:39]
  assign pes_38_io_cfg_data = cfgRegs_26[31:0]; // @[CGRA.scala 673:39]
  assign pes_38_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_38_io_in_0 = gibs_50_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_38_io_in_1 = gibs_51_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_38_io_in_2 = gibs_54_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_38_io_in_3 = gibs_55_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_38_io_in_4 = gibs_50_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_38_io_in_5 = gibs_51_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_38_io_in_6 = gibs_54_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_38_io_in_7 = gibs_55_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_39_clock = clock;
  assign pes_39_reset = reset;
  assign pes_39_io_cfg_en = cfgRegs_28[46]; // @[CGRA.scala 671:37]
  assign pes_39_io_cfg_addr = cfgRegs_28[45:32]; // @[CGRA.scala 672:39]
  assign pes_39_io_cfg_data = cfgRegs_28[31:0]; // @[CGRA.scala 673:39]
  assign pes_39_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_39_io_in_0 = gibs_52_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_39_io_in_1 = gibs_53_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_39_io_in_2 = gibs_56_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_39_io_in_3 = gibs_57_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_39_io_in_4 = gibs_52_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_39_io_in_5 = gibs_53_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_39_io_in_6 = gibs_56_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_39_io_in_7 = gibs_57_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_40_clock = clock;
  assign pes_40_reset = reset;
  assign pes_40_io_cfg_en = cfgRegs_28[46]; // @[CGRA.scala 671:37]
  assign pes_40_io_cfg_addr = cfgRegs_28[45:32]; // @[CGRA.scala 672:39]
  assign pes_40_io_cfg_data = cfgRegs_28[31:0]; // @[CGRA.scala 673:39]
  assign pes_40_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_40_io_in_0 = gibs_53_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_40_io_in_1 = gibs_54_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_40_io_in_2 = gibs_57_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_40_io_in_3 = gibs_58_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_40_io_in_4 = gibs_53_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_40_io_in_5 = gibs_54_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_40_io_in_6 = gibs_57_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_40_io_in_7 = gibs_58_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_41_clock = clock;
  assign pes_41_reset = reset;
  assign pes_41_io_cfg_en = cfgRegs_28[46]; // @[CGRA.scala 671:37]
  assign pes_41_io_cfg_addr = cfgRegs_28[45:32]; // @[CGRA.scala 672:39]
  assign pes_41_io_cfg_data = cfgRegs_28[31:0]; // @[CGRA.scala 673:39]
  assign pes_41_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_41_io_in_0 = gibs_54_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_41_io_in_1 = gibs_55_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_41_io_in_2 = gibs_58_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_41_io_in_3 = gibs_59_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_41_io_in_4 = gibs_54_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_41_io_in_5 = gibs_55_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_41_io_in_6 = gibs_58_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_41_io_in_7 = gibs_59_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_42_clock = clock;
  assign pes_42_reset = reset;
  assign pes_42_io_cfg_en = cfgRegs_30[46]; // @[CGRA.scala 671:37]
  assign pes_42_io_cfg_addr = cfgRegs_30[45:32]; // @[CGRA.scala 672:39]
  assign pes_42_io_cfg_data = cfgRegs_30[31:0]; // @[CGRA.scala 673:39]
  assign pes_42_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_42_io_in_0 = gibs_56_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_42_io_in_1 = gibs_57_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_42_io_in_2 = gibs_60_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_42_io_in_3 = gibs_61_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_42_io_in_4 = gibs_56_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_42_io_in_5 = gibs_57_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_42_io_in_6 = gibs_60_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_42_io_in_7 = gibs_61_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_43_clock = clock;
  assign pes_43_reset = reset;
  assign pes_43_io_cfg_en = cfgRegs_30[46]; // @[CGRA.scala 671:37]
  assign pes_43_io_cfg_addr = cfgRegs_30[45:32]; // @[CGRA.scala 672:39]
  assign pes_43_io_cfg_data = cfgRegs_30[31:0]; // @[CGRA.scala 673:39]
  assign pes_43_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_43_io_in_0 = gibs_57_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_43_io_in_1 = gibs_58_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_43_io_in_2 = gibs_61_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_43_io_in_3 = gibs_62_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_43_io_in_4 = gibs_57_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_43_io_in_5 = gibs_58_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_43_io_in_6 = gibs_61_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_43_io_in_7 = gibs_62_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_44_clock = clock;
  assign pes_44_reset = reset;
  assign pes_44_io_cfg_en = cfgRegs_30[46]; // @[CGRA.scala 671:37]
  assign pes_44_io_cfg_addr = cfgRegs_30[45:32]; // @[CGRA.scala 672:39]
  assign pes_44_io_cfg_data = cfgRegs_30[31:0]; // @[CGRA.scala 673:39]
  assign pes_44_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_44_io_in_0 = gibs_58_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_44_io_in_1 = gibs_59_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_44_io_in_2 = gibs_62_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_44_io_in_3 = gibs_63_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_44_io_in_4 = gibs_58_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_44_io_in_5 = gibs_59_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_44_io_in_6 = gibs_62_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_44_io_in_7 = gibs_63_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_45_clock = clock;
  assign pes_45_reset = reset;
  assign pes_45_io_cfg_en = cfgRegs_32[46]; // @[CGRA.scala 671:37]
  assign pes_45_io_cfg_addr = cfgRegs_32[45:32]; // @[CGRA.scala 672:39]
  assign pes_45_io_cfg_data = cfgRegs_32[31:0]; // @[CGRA.scala 673:39]
  assign pes_45_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_45_io_in_0 = gibs_60_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_45_io_in_1 = gibs_61_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_45_io_in_2 = gibs_64_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_45_io_in_3 = gibs_65_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_45_io_in_4 = gibs_60_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_45_io_in_5 = gibs_61_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_45_io_in_6 = gibs_64_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_45_io_in_7 = gibs_65_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_46_clock = clock;
  assign pes_46_reset = reset;
  assign pes_46_io_cfg_en = cfgRegs_32[46]; // @[CGRA.scala 671:37]
  assign pes_46_io_cfg_addr = cfgRegs_32[45:32]; // @[CGRA.scala 672:39]
  assign pes_46_io_cfg_data = cfgRegs_32[31:0]; // @[CGRA.scala 673:39]
  assign pes_46_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_46_io_in_0 = gibs_61_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_46_io_in_1 = gibs_62_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_46_io_in_2 = gibs_65_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_46_io_in_3 = gibs_66_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_46_io_in_4 = gibs_61_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_46_io_in_5 = gibs_62_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_46_io_in_6 = gibs_65_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_46_io_in_7 = gibs_66_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_47_clock = clock;
  assign pes_47_reset = reset;
  assign pes_47_io_cfg_en = cfgRegs_32[46]; // @[CGRA.scala 671:37]
  assign pes_47_io_cfg_addr = cfgRegs_32[45:32]; // @[CGRA.scala 672:39]
  assign pes_47_io_cfg_data = cfgRegs_32[31:0]; // @[CGRA.scala 673:39]
  assign pes_47_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_47_io_in_0 = gibs_62_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_47_io_in_1 = gibs_63_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_47_io_in_2 = gibs_66_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_47_io_in_3 = gibs_67_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_47_io_in_4 = gibs_62_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_47_io_in_5 = gibs_63_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_47_io_in_6 = gibs_66_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_47_io_in_7 = gibs_67_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_48_clock = clock;
  assign pes_48_reset = reset;
  assign pes_48_io_cfg_en = cfgRegs_34[46]; // @[CGRA.scala 671:37]
  assign pes_48_io_cfg_addr = cfgRegs_34[45:32]; // @[CGRA.scala 672:39]
  assign pes_48_io_cfg_data = cfgRegs_34[31:0]; // @[CGRA.scala 673:39]
  assign pes_48_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_48_io_in_0 = gibs_64_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_48_io_in_1 = gibs_65_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_48_io_in_2 = gibs_68_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_48_io_in_3 = gibs_69_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_48_io_in_4 = gibs_64_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_48_io_in_5 = gibs_65_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_48_io_in_6 = gibs_68_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_48_io_in_7 = gibs_69_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_49_clock = clock;
  assign pes_49_reset = reset;
  assign pes_49_io_cfg_en = cfgRegs_34[46]; // @[CGRA.scala 671:37]
  assign pes_49_io_cfg_addr = cfgRegs_34[45:32]; // @[CGRA.scala 672:39]
  assign pes_49_io_cfg_data = cfgRegs_34[31:0]; // @[CGRA.scala 673:39]
  assign pes_49_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_49_io_in_0 = gibs_65_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_49_io_in_1 = gibs_66_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_49_io_in_2 = gibs_69_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_49_io_in_3 = gibs_70_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_49_io_in_4 = gibs_65_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_49_io_in_5 = gibs_66_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_49_io_in_6 = gibs_69_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_49_io_in_7 = gibs_70_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_50_clock = clock;
  assign pes_50_reset = reset;
  assign pes_50_io_cfg_en = cfgRegs_34[46]; // @[CGRA.scala 671:37]
  assign pes_50_io_cfg_addr = cfgRegs_34[45:32]; // @[CGRA.scala 672:39]
  assign pes_50_io_cfg_data = cfgRegs_34[31:0]; // @[CGRA.scala 673:39]
  assign pes_50_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_50_io_in_0 = gibs_66_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_50_io_in_1 = gibs_67_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_50_io_in_2 = gibs_70_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_50_io_in_3 = gibs_71_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_50_io_in_4 = gibs_66_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_50_io_in_5 = gibs_67_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_50_io_in_6 = gibs_70_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_50_io_in_7 = gibs_71_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_51_clock = clock;
  assign pes_51_reset = reset;
  assign pes_51_io_cfg_en = cfgRegs_36[46]; // @[CGRA.scala 671:37]
  assign pes_51_io_cfg_addr = cfgRegs_36[45:32]; // @[CGRA.scala 672:39]
  assign pes_51_io_cfg_data = cfgRegs_36[31:0]; // @[CGRA.scala 673:39]
  assign pes_51_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_51_io_in_0 = gibs_68_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_51_io_in_1 = gibs_69_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_51_io_in_2 = gibs_72_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_51_io_in_3 = gibs_73_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_51_io_in_4 = gibs_68_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_51_io_in_5 = gibs_69_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_51_io_in_6 = gibs_72_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_51_io_in_7 = gibs_73_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_52_clock = clock;
  assign pes_52_reset = reset;
  assign pes_52_io_cfg_en = cfgRegs_36[46]; // @[CGRA.scala 671:37]
  assign pes_52_io_cfg_addr = cfgRegs_36[45:32]; // @[CGRA.scala 672:39]
  assign pes_52_io_cfg_data = cfgRegs_36[31:0]; // @[CGRA.scala 673:39]
  assign pes_52_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_52_io_in_0 = gibs_69_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_52_io_in_1 = gibs_70_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_52_io_in_2 = gibs_73_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_52_io_in_3 = gibs_74_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_52_io_in_4 = gibs_69_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_52_io_in_5 = gibs_70_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_52_io_in_6 = gibs_73_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_52_io_in_7 = gibs_74_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_53_clock = clock;
  assign pes_53_reset = reset;
  assign pes_53_io_cfg_en = cfgRegs_36[46]; // @[CGRA.scala 671:37]
  assign pes_53_io_cfg_addr = cfgRegs_36[45:32]; // @[CGRA.scala 672:39]
  assign pes_53_io_cfg_data = cfgRegs_36[31:0]; // @[CGRA.scala 673:39]
  assign pes_53_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_53_io_in_0 = gibs_70_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_53_io_in_1 = gibs_71_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_53_io_in_2 = gibs_74_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_53_io_in_3 = gibs_75_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_53_io_in_4 = gibs_70_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_53_io_in_5 = gibs_71_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_53_io_in_6 = gibs_74_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_53_io_in_7 = gibs_75_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_54_clock = clock;
  assign pes_54_reset = reset;
  assign pes_54_io_cfg_en = cfgRegs_38[46]; // @[CGRA.scala 671:37]
  assign pes_54_io_cfg_addr = cfgRegs_38[45:32]; // @[CGRA.scala 672:39]
  assign pes_54_io_cfg_data = cfgRegs_38[31:0]; // @[CGRA.scala 673:39]
  assign pes_54_io_en = io_en_1; // @[CGRA.scala 476:27]
  assign pes_54_io_in_0 = gibs_72_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_54_io_in_1 = gibs_73_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_54_io_in_2 = gibs_76_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_54_io_in_3 = gibs_77_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_54_io_in_4 = gibs_72_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_54_io_in_5 = gibs_73_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_54_io_in_6 = gibs_76_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_54_io_in_7 = gibs_77_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_55_clock = clock;
  assign pes_55_reset = reset;
  assign pes_55_io_cfg_en = cfgRegs_38[46]; // @[CGRA.scala 671:37]
  assign pes_55_io_cfg_addr = cfgRegs_38[45:32]; // @[CGRA.scala 672:39]
  assign pes_55_io_cfg_data = cfgRegs_38[31:0]; // @[CGRA.scala 673:39]
  assign pes_55_io_en = io_en_2; // @[CGRA.scala 476:27]
  assign pes_55_io_in_0 = gibs_73_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_55_io_in_1 = gibs_74_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_55_io_in_2 = gibs_77_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_55_io_in_3 = gibs_78_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_55_io_in_4 = gibs_73_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_55_io_in_5 = gibs_74_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_55_io_in_6 = gibs_77_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_55_io_in_7 = gibs_78_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign pes_56_clock = clock;
  assign pes_56_reset = reset;
  assign pes_56_io_cfg_en = cfgRegs_38[46]; // @[CGRA.scala 671:37]
  assign pes_56_io_cfg_addr = cfgRegs_38[45:32]; // @[CGRA.scala 672:39]
  assign pes_56_io_cfg_data = cfgRegs_38[31:0]; // @[CGRA.scala 673:39]
  assign pes_56_io_en = io_en_3; // @[CGRA.scala 476:27]
  assign pes_56_io_in_0 = gibs_74_io_ipinSE_0; // @[CGRA.scala 479:14]
  assign pes_56_io_in_1 = gibs_75_io_ipinSW_0; // @[CGRA.scala 483:14]
  assign pes_56_io_in_2 = gibs_78_io_ipinNE_0; // @[CGRA.scala 487:14]
  assign pes_56_io_in_3 = gibs_79_io_ipinNW_0; // @[CGRA.scala 491:14]
  assign pes_56_io_in_4 = gibs_74_io_ipinSE_1; // @[CGRA.scala 479:14]
  assign pes_56_io_in_5 = gibs_75_io_ipinSW_1; // @[CGRA.scala 483:14]
  assign pes_56_io_in_6 = gibs_78_io_ipinNE_1; // @[CGRA.scala 487:14]
  assign pes_56_io_in_7 = gibs_79_io_ipinNW_1; // @[CGRA.scala 491:14]
  assign gibs_0_clock = clock;
  assign gibs_0_reset = reset;
  assign gibs_0_io_cfg_en = cfgRegs_1[46]; // @[CGRA.scala 667:42]
  assign gibs_0_io_cfg_addr = cfgRegs_1[45:32]; // @[CGRA.scala 668:44]
  assign gibs_0_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 669:44]
  assign gibs_0_io_opinNE_0 = ibs_0_io_out_0; // @[CGRA.scala 420:35]
  assign gibs_0_io_opinSE_0 = pes_0_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_0_io_opinSW_0 = lsus_0_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_0_io_itrackE_0 = gibs_1_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_0_io_itrackS_0 = gibs_4_io_otrackN_0; // @[CGRA.scala 521:16]
  assign gibs_1_clock = clock;
  assign gibs_1_reset = reset;
  assign gibs_1_io_cfg_en = cfgRegs_1[46]; // @[CGRA.scala 667:42]
  assign gibs_1_io_cfg_addr = cfgRegs_1[45:32]; // @[CGRA.scala 668:44]
  assign gibs_1_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 669:44]
  assign gibs_1_io_opinNW_0 = ibs_0_io_out_0; // @[CGRA.scala 421:37]
  assign gibs_1_io_opinNE_0 = ibs_1_io_out_0; // @[CGRA.scala 420:35]
  assign gibs_1_io_opinSE_0 = pes_1_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_1_io_opinSW_0 = pes_0_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_1_io_itrackW_0 = gibs_0_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_1_io_itrackE_0 = gibs_2_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_1_io_itrackS_0 = gibs_5_io_otrackN_0; // @[CGRA.scala 521:16]
  assign gibs_2_clock = clock;
  assign gibs_2_reset = reset;
  assign gibs_2_io_cfg_en = cfgRegs_1[46]; // @[CGRA.scala 667:42]
  assign gibs_2_io_cfg_addr = cfgRegs_1[45:32]; // @[CGRA.scala 668:44]
  assign gibs_2_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 669:44]
  assign gibs_2_io_opinNW_0 = ibs_1_io_out_0; // @[CGRA.scala 421:37]
  assign gibs_2_io_opinNE_0 = ibs_2_io_out_0; // @[CGRA.scala 420:35]
  assign gibs_2_io_opinSE_0 = pes_2_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_2_io_opinSW_0 = pes_1_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_2_io_itrackW_0 = gibs_1_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_2_io_itrackE_0 = gibs_3_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_2_io_itrackS_0 = gibs_6_io_otrackN_0; // @[CGRA.scala 521:16]
  assign gibs_3_clock = clock;
  assign gibs_3_reset = reset;
  assign gibs_3_io_cfg_en = cfgRegs_1[46]; // @[CGRA.scala 667:42]
  assign gibs_3_io_cfg_addr = cfgRegs_1[45:32]; // @[CGRA.scala 668:44]
  assign gibs_3_io_cfg_data = cfgRegs_1[31:0]; // @[CGRA.scala 669:44]
  assign gibs_3_io_opinNW_0 = ibs_2_io_out_0; // @[CGRA.scala 421:37]
  assign gibs_3_io_opinSE_0 = lsus_1_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_3_io_opinSW_0 = pes_2_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_3_io_itrackW_0 = gibs_2_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_3_io_itrackS_0 = gibs_7_io_otrackN_0; // @[CGRA.scala 521:16]
  assign gibs_4_clock = clock;
  assign gibs_4_reset = reset;
  assign gibs_4_io_cfg_en = cfgRegs_3[46]; // @[CGRA.scala 667:42]
  assign gibs_4_io_cfg_addr = cfgRegs_3[45:32]; // @[CGRA.scala 668:44]
  assign gibs_4_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 669:44]
  assign gibs_4_io_opinNW_0 = lsus_0_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_4_io_opinNE_0 = pes_0_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_4_io_opinSE_0 = pes_3_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_4_io_opinSW_0 = lsus_2_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_4_io_itrackN_0 = gibs_0_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_4_io_itrackE_0 = gibs_5_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_4_io_itrackS_0 = gibs_8_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_5_clock = clock;
  assign gibs_5_reset = reset;
  assign gibs_5_io_cfg_en = cfgRegs_3[46]; // @[CGRA.scala 667:42]
  assign gibs_5_io_cfg_addr = cfgRegs_3[45:32]; // @[CGRA.scala 668:44]
  assign gibs_5_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 669:44]
  assign gibs_5_io_opinNW_0 = pes_0_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_5_io_opinNE_0 = pes_1_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_5_io_opinSE_0 = pes_4_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_5_io_opinSW_0 = pes_3_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_5_io_itrackW_0 = gibs_4_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_5_io_itrackN_0 = gibs_1_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_5_io_itrackE_0 = gibs_6_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_5_io_itrackS_0 = gibs_9_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_6_clock = clock;
  assign gibs_6_reset = reset;
  assign gibs_6_io_cfg_en = cfgRegs_3[46]; // @[CGRA.scala 667:42]
  assign gibs_6_io_cfg_addr = cfgRegs_3[45:32]; // @[CGRA.scala 668:44]
  assign gibs_6_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 669:44]
  assign gibs_6_io_opinNW_0 = pes_1_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_6_io_opinNE_0 = pes_2_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_6_io_opinSE_0 = pes_5_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_6_io_opinSW_0 = pes_4_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_6_io_itrackW_0 = gibs_5_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_6_io_itrackN_0 = gibs_2_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_6_io_itrackE_0 = gibs_7_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_6_io_itrackS_0 = gibs_10_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_7_clock = clock;
  assign gibs_7_reset = reset;
  assign gibs_7_io_cfg_en = cfgRegs_3[46]; // @[CGRA.scala 667:42]
  assign gibs_7_io_cfg_addr = cfgRegs_3[45:32]; // @[CGRA.scala 668:44]
  assign gibs_7_io_cfg_data = cfgRegs_3[31:0]; // @[CGRA.scala 669:44]
  assign gibs_7_io_opinNW_0 = pes_2_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_7_io_opinNE_0 = lsus_1_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_7_io_opinSE_0 = lsus_3_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_7_io_opinSW_0 = pes_5_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_7_io_itrackW_0 = gibs_6_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_7_io_itrackN_0 = gibs_3_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_7_io_itrackS_0 = gibs_11_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_8_clock = clock;
  assign gibs_8_reset = reset;
  assign gibs_8_io_cfg_en = cfgRegs_5[46]; // @[CGRA.scala 667:42]
  assign gibs_8_io_cfg_addr = cfgRegs_5[45:32]; // @[CGRA.scala 668:44]
  assign gibs_8_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 669:44]
  assign gibs_8_io_opinNW_0 = lsus_2_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_8_io_opinNE_0 = pes_3_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_8_io_opinSE_0 = pes_6_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_8_io_opinSW_0 = lsus_4_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_8_io_itrackN_0 = gibs_4_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_8_io_itrackE_0 = gibs_9_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_8_io_itrackS_0 = gibs_12_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_9_clock = clock;
  assign gibs_9_reset = reset;
  assign gibs_9_io_cfg_en = cfgRegs_5[46]; // @[CGRA.scala 667:42]
  assign gibs_9_io_cfg_addr = cfgRegs_5[45:32]; // @[CGRA.scala 668:44]
  assign gibs_9_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 669:44]
  assign gibs_9_io_opinNW_0 = pes_3_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_9_io_opinNE_0 = pes_4_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_9_io_opinSE_0 = pes_7_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_9_io_opinSW_0 = pes_6_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_9_io_itrackW_0 = gibs_8_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_9_io_itrackN_0 = gibs_5_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_9_io_itrackE_0 = gibs_10_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_9_io_itrackS_0 = gibs_13_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_10_clock = clock;
  assign gibs_10_reset = reset;
  assign gibs_10_io_cfg_en = cfgRegs_5[46]; // @[CGRA.scala 667:42]
  assign gibs_10_io_cfg_addr = cfgRegs_5[45:32]; // @[CGRA.scala 668:44]
  assign gibs_10_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 669:44]
  assign gibs_10_io_opinNW_0 = pes_4_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_10_io_opinNE_0 = pes_5_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_10_io_opinSE_0 = pes_8_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_10_io_opinSW_0 = pes_7_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_10_io_itrackW_0 = gibs_9_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_10_io_itrackN_0 = gibs_6_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_10_io_itrackE_0 = gibs_11_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_10_io_itrackS_0 = gibs_14_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_11_clock = clock;
  assign gibs_11_reset = reset;
  assign gibs_11_io_cfg_en = cfgRegs_5[46]; // @[CGRA.scala 667:42]
  assign gibs_11_io_cfg_addr = cfgRegs_5[45:32]; // @[CGRA.scala 668:44]
  assign gibs_11_io_cfg_data = cfgRegs_5[31:0]; // @[CGRA.scala 669:44]
  assign gibs_11_io_opinNW_0 = pes_5_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_11_io_opinNE_0 = lsus_3_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_11_io_opinSE_0 = lsus_5_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_11_io_opinSW_0 = pes_8_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_11_io_itrackW_0 = gibs_10_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_11_io_itrackN_0 = gibs_7_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_11_io_itrackS_0 = gibs_15_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_12_clock = clock;
  assign gibs_12_reset = reset;
  assign gibs_12_io_cfg_en = cfgRegs_7[46]; // @[CGRA.scala 667:42]
  assign gibs_12_io_cfg_addr = cfgRegs_7[45:32]; // @[CGRA.scala 668:44]
  assign gibs_12_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 669:44]
  assign gibs_12_io_opinNW_0 = lsus_4_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_12_io_opinNE_0 = pes_6_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_12_io_opinSE_0 = pes_9_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_12_io_opinSW_0 = lsus_6_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_12_io_itrackN_0 = gibs_8_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_12_io_itrackE_0 = gibs_13_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_12_io_itrackS_0 = gibs_16_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_13_clock = clock;
  assign gibs_13_reset = reset;
  assign gibs_13_io_cfg_en = cfgRegs_7[46]; // @[CGRA.scala 667:42]
  assign gibs_13_io_cfg_addr = cfgRegs_7[45:32]; // @[CGRA.scala 668:44]
  assign gibs_13_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 669:44]
  assign gibs_13_io_opinNW_0 = pes_6_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_13_io_opinNE_0 = pes_7_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_13_io_opinSE_0 = pes_10_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_13_io_opinSW_0 = pes_9_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_13_io_itrackW_0 = gibs_12_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_13_io_itrackN_0 = gibs_9_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_13_io_itrackE_0 = gibs_14_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_13_io_itrackS_0 = gibs_17_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_14_clock = clock;
  assign gibs_14_reset = reset;
  assign gibs_14_io_cfg_en = cfgRegs_7[46]; // @[CGRA.scala 667:42]
  assign gibs_14_io_cfg_addr = cfgRegs_7[45:32]; // @[CGRA.scala 668:44]
  assign gibs_14_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 669:44]
  assign gibs_14_io_opinNW_0 = pes_7_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_14_io_opinNE_0 = pes_8_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_14_io_opinSE_0 = pes_11_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_14_io_opinSW_0 = pes_10_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_14_io_itrackW_0 = gibs_13_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_14_io_itrackN_0 = gibs_10_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_14_io_itrackE_0 = gibs_15_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_14_io_itrackS_0 = gibs_18_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_15_clock = clock;
  assign gibs_15_reset = reset;
  assign gibs_15_io_cfg_en = cfgRegs_7[46]; // @[CGRA.scala 667:42]
  assign gibs_15_io_cfg_addr = cfgRegs_7[45:32]; // @[CGRA.scala 668:44]
  assign gibs_15_io_cfg_data = cfgRegs_7[31:0]; // @[CGRA.scala 669:44]
  assign gibs_15_io_opinNW_0 = pes_8_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_15_io_opinNE_0 = lsus_5_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_15_io_opinSE_0 = lsus_7_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_15_io_opinSW_0 = pes_11_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_15_io_itrackW_0 = gibs_14_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_15_io_itrackN_0 = gibs_11_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_15_io_itrackS_0 = gibs_19_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_16_clock = clock;
  assign gibs_16_reset = reset;
  assign gibs_16_io_cfg_en = cfgRegs_9[46]; // @[CGRA.scala 667:42]
  assign gibs_16_io_cfg_addr = cfgRegs_9[45:32]; // @[CGRA.scala 668:44]
  assign gibs_16_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 669:44]
  assign gibs_16_io_opinNW_0 = lsus_6_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_16_io_opinNE_0 = pes_9_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_16_io_opinSE_0 = pes_12_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_16_io_opinSW_0 = lsus_8_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_16_io_itrackN_0 = gibs_12_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_16_io_itrackE_0 = gibs_17_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_16_io_itrackS_0 = gibs_20_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_17_clock = clock;
  assign gibs_17_reset = reset;
  assign gibs_17_io_cfg_en = cfgRegs_9[46]; // @[CGRA.scala 667:42]
  assign gibs_17_io_cfg_addr = cfgRegs_9[45:32]; // @[CGRA.scala 668:44]
  assign gibs_17_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 669:44]
  assign gibs_17_io_opinNW_0 = pes_9_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_17_io_opinNE_0 = pes_10_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_17_io_opinSE_0 = pes_13_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_17_io_opinSW_0 = pes_12_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_17_io_itrackW_0 = gibs_16_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_17_io_itrackN_0 = gibs_13_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_17_io_itrackE_0 = gibs_18_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_17_io_itrackS_0 = gibs_21_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_18_clock = clock;
  assign gibs_18_reset = reset;
  assign gibs_18_io_cfg_en = cfgRegs_9[46]; // @[CGRA.scala 667:42]
  assign gibs_18_io_cfg_addr = cfgRegs_9[45:32]; // @[CGRA.scala 668:44]
  assign gibs_18_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 669:44]
  assign gibs_18_io_opinNW_0 = pes_10_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_18_io_opinNE_0 = pes_11_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_18_io_opinSE_0 = pes_14_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_18_io_opinSW_0 = pes_13_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_18_io_itrackW_0 = gibs_17_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_18_io_itrackN_0 = gibs_14_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_18_io_itrackE_0 = gibs_19_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_18_io_itrackS_0 = gibs_22_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_19_clock = clock;
  assign gibs_19_reset = reset;
  assign gibs_19_io_cfg_en = cfgRegs_9[46]; // @[CGRA.scala 667:42]
  assign gibs_19_io_cfg_addr = cfgRegs_9[45:32]; // @[CGRA.scala 668:44]
  assign gibs_19_io_cfg_data = cfgRegs_9[31:0]; // @[CGRA.scala 669:44]
  assign gibs_19_io_opinNW_0 = pes_11_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_19_io_opinNE_0 = lsus_7_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_19_io_opinSE_0 = lsus_9_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_19_io_opinSW_0 = pes_14_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_19_io_itrackW_0 = gibs_18_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_19_io_itrackN_0 = gibs_15_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_19_io_itrackS_0 = gibs_23_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_20_clock = clock;
  assign gibs_20_reset = reset;
  assign gibs_20_io_cfg_en = cfgRegs_11[46]; // @[CGRA.scala 667:42]
  assign gibs_20_io_cfg_addr = cfgRegs_11[45:32]; // @[CGRA.scala 668:44]
  assign gibs_20_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 669:44]
  assign gibs_20_io_opinNW_0 = lsus_8_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_20_io_opinNE_0 = pes_12_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_20_io_opinSE_0 = pes_15_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_20_io_opinSW_0 = lsus_10_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_20_io_itrackN_0 = gibs_16_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_20_io_itrackE_0 = gibs_21_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_20_io_itrackS_0 = gibs_24_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_21_clock = clock;
  assign gibs_21_reset = reset;
  assign gibs_21_io_cfg_en = cfgRegs_11[46]; // @[CGRA.scala 667:42]
  assign gibs_21_io_cfg_addr = cfgRegs_11[45:32]; // @[CGRA.scala 668:44]
  assign gibs_21_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 669:44]
  assign gibs_21_io_opinNW_0 = pes_12_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_21_io_opinNE_0 = pes_13_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_21_io_opinSE_0 = pes_16_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_21_io_opinSW_0 = pes_15_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_21_io_itrackW_0 = gibs_20_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_21_io_itrackN_0 = gibs_17_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_21_io_itrackE_0 = gibs_22_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_21_io_itrackS_0 = gibs_25_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_22_clock = clock;
  assign gibs_22_reset = reset;
  assign gibs_22_io_cfg_en = cfgRegs_11[46]; // @[CGRA.scala 667:42]
  assign gibs_22_io_cfg_addr = cfgRegs_11[45:32]; // @[CGRA.scala 668:44]
  assign gibs_22_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 669:44]
  assign gibs_22_io_opinNW_0 = pes_13_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_22_io_opinNE_0 = pes_14_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_22_io_opinSE_0 = pes_17_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_22_io_opinSW_0 = pes_16_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_22_io_itrackW_0 = gibs_21_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_22_io_itrackN_0 = gibs_18_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_22_io_itrackE_0 = gibs_23_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_22_io_itrackS_0 = gibs_26_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_23_clock = clock;
  assign gibs_23_reset = reset;
  assign gibs_23_io_cfg_en = cfgRegs_11[46]; // @[CGRA.scala 667:42]
  assign gibs_23_io_cfg_addr = cfgRegs_11[45:32]; // @[CGRA.scala 668:44]
  assign gibs_23_io_cfg_data = cfgRegs_11[31:0]; // @[CGRA.scala 669:44]
  assign gibs_23_io_opinNW_0 = pes_14_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_23_io_opinNE_0 = lsus_9_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_23_io_opinSE_0 = lsus_11_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_23_io_opinSW_0 = pes_17_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_23_io_itrackW_0 = gibs_22_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_23_io_itrackN_0 = gibs_19_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_23_io_itrackS_0 = gibs_27_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_24_clock = clock;
  assign gibs_24_reset = reset;
  assign gibs_24_io_cfg_en = cfgRegs_13[46]; // @[CGRA.scala 667:42]
  assign gibs_24_io_cfg_addr = cfgRegs_13[45:32]; // @[CGRA.scala 668:44]
  assign gibs_24_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 669:44]
  assign gibs_24_io_opinNW_0 = lsus_10_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_24_io_opinNE_0 = pes_15_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_24_io_opinSE_0 = pes_18_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_24_io_opinSW_0 = lsus_12_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_24_io_itrackN_0 = gibs_20_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_24_io_itrackE_0 = gibs_25_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_24_io_itrackS_0 = gibs_28_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_25_clock = clock;
  assign gibs_25_reset = reset;
  assign gibs_25_io_cfg_en = cfgRegs_13[46]; // @[CGRA.scala 667:42]
  assign gibs_25_io_cfg_addr = cfgRegs_13[45:32]; // @[CGRA.scala 668:44]
  assign gibs_25_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 669:44]
  assign gibs_25_io_opinNW_0 = pes_15_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_25_io_opinNE_0 = pes_16_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_25_io_opinSE_0 = pes_19_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_25_io_opinSW_0 = pes_18_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_25_io_itrackW_0 = gibs_24_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_25_io_itrackN_0 = gibs_21_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_25_io_itrackE_0 = gibs_26_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_25_io_itrackS_0 = gibs_29_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_26_clock = clock;
  assign gibs_26_reset = reset;
  assign gibs_26_io_cfg_en = cfgRegs_13[46]; // @[CGRA.scala 667:42]
  assign gibs_26_io_cfg_addr = cfgRegs_13[45:32]; // @[CGRA.scala 668:44]
  assign gibs_26_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 669:44]
  assign gibs_26_io_opinNW_0 = pes_16_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_26_io_opinNE_0 = pes_17_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_26_io_opinSE_0 = pes_20_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_26_io_opinSW_0 = pes_19_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_26_io_itrackW_0 = gibs_25_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_26_io_itrackN_0 = gibs_22_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_26_io_itrackE_0 = gibs_27_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_26_io_itrackS_0 = gibs_30_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_27_clock = clock;
  assign gibs_27_reset = reset;
  assign gibs_27_io_cfg_en = cfgRegs_13[46]; // @[CGRA.scala 667:42]
  assign gibs_27_io_cfg_addr = cfgRegs_13[45:32]; // @[CGRA.scala 668:44]
  assign gibs_27_io_cfg_data = cfgRegs_13[31:0]; // @[CGRA.scala 669:44]
  assign gibs_27_io_opinNW_0 = pes_17_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_27_io_opinNE_0 = lsus_11_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_27_io_opinSE_0 = lsus_13_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_27_io_opinSW_0 = pes_20_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_27_io_itrackW_0 = gibs_26_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_27_io_itrackN_0 = gibs_23_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_27_io_itrackS_0 = gibs_31_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_28_clock = clock;
  assign gibs_28_reset = reset;
  assign gibs_28_io_cfg_en = cfgRegs_15[46]; // @[CGRA.scala 667:42]
  assign gibs_28_io_cfg_addr = cfgRegs_15[45:32]; // @[CGRA.scala 668:44]
  assign gibs_28_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 669:44]
  assign gibs_28_io_opinNW_0 = lsus_12_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_28_io_opinNE_0 = pes_18_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_28_io_opinSE_0 = pes_21_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_28_io_opinSW_0 = lsus_14_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_28_io_itrackN_0 = gibs_24_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_28_io_itrackE_0 = gibs_29_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_28_io_itrackS_0 = gibs_32_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_29_clock = clock;
  assign gibs_29_reset = reset;
  assign gibs_29_io_cfg_en = cfgRegs_15[46]; // @[CGRA.scala 667:42]
  assign gibs_29_io_cfg_addr = cfgRegs_15[45:32]; // @[CGRA.scala 668:44]
  assign gibs_29_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 669:44]
  assign gibs_29_io_opinNW_0 = pes_18_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_29_io_opinNE_0 = pes_19_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_29_io_opinSE_0 = pes_22_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_29_io_opinSW_0 = pes_21_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_29_io_itrackW_0 = gibs_28_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_29_io_itrackN_0 = gibs_25_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_29_io_itrackE_0 = gibs_30_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_29_io_itrackS_0 = gibs_33_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_30_clock = clock;
  assign gibs_30_reset = reset;
  assign gibs_30_io_cfg_en = cfgRegs_15[46]; // @[CGRA.scala 667:42]
  assign gibs_30_io_cfg_addr = cfgRegs_15[45:32]; // @[CGRA.scala 668:44]
  assign gibs_30_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 669:44]
  assign gibs_30_io_opinNW_0 = pes_19_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_30_io_opinNE_0 = pes_20_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_30_io_opinSE_0 = pes_23_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_30_io_opinSW_0 = pes_22_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_30_io_itrackW_0 = gibs_29_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_30_io_itrackN_0 = gibs_26_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_30_io_itrackE_0 = gibs_31_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_30_io_itrackS_0 = gibs_34_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_31_clock = clock;
  assign gibs_31_reset = reset;
  assign gibs_31_io_cfg_en = cfgRegs_15[46]; // @[CGRA.scala 667:42]
  assign gibs_31_io_cfg_addr = cfgRegs_15[45:32]; // @[CGRA.scala 668:44]
  assign gibs_31_io_cfg_data = cfgRegs_15[31:0]; // @[CGRA.scala 669:44]
  assign gibs_31_io_opinNW_0 = pes_20_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_31_io_opinNE_0 = lsus_13_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_31_io_opinSE_0 = lsus_15_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_31_io_opinSW_0 = pes_23_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_31_io_itrackW_0 = gibs_30_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_31_io_itrackN_0 = gibs_27_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_31_io_itrackS_0 = gibs_35_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_32_clock = clock;
  assign gibs_32_reset = reset;
  assign gibs_32_io_cfg_en = cfgRegs_17[46]; // @[CGRA.scala 667:42]
  assign gibs_32_io_cfg_addr = cfgRegs_17[45:32]; // @[CGRA.scala 668:44]
  assign gibs_32_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 669:44]
  assign gibs_32_io_opinNW_0 = lsus_14_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_32_io_opinNE_0 = pes_21_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_32_io_opinSE_0 = pes_24_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_32_io_opinSW_0 = lsus_16_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_32_io_itrackN_0 = gibs_28_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_32_io_itrackE_0 = gibs_33_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_32_io_itrackS_0 = gibs_36_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_33_clock = clock;
  assign gibs_33_reset = reset;
  assign gibs_33_io_cfg_en = cfgRegs_17[46]; // @[CGRA.scala 667:42]
  assign gibs_33_io_cfg_addr = cfgRegs_17[45:32]; // @[CGRA.scala 668:44]
  assign gibs_33_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 669:44]
  assign gibs_33_io_opinNW_0 = pes_21_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_33_io_opinNE_0 = pes_22_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_33_io_opinSE_0 = pes_25_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_33_io_opinSW_0 = pes_24_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_33_io_itrackW_0 = gibs_32_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_33_io_itrackN_0 = gibs_29_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_33_io_itrackE_0 = gibs_34_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_33_io_itrackS_0 = gibs_37_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_34_clock = clock;
  assign gibs_34_reset = reset;
  assign gibs_34_io_cfg_en = cfgRegs_17[46]; // @[CGRA.scala 667:42]
  assign gibs_34_io_cfg_addr = cfgRegs_17[45:32]; // @[CGRA.scala 668:44]
  assign gibs_34_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 669:44]
  assign gibs_34_io_opinNW_0 = pes_22_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_34_io_opinNE_0 = pes_23_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_34_io_opinSE_0 = pes_26_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_34_io_opinSW_0 = pes_25_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_34_io_itrackW_0 = gibs_33_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_34_io_itrackN_0 = gibs_30_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_34_io_itrackE_0 = gibs_35_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_34_io_itrackS_0 = gibs_38_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_35_clock = clock;
  assign gibs_35_reset = reset;
  assign gibs_35_io_cfg_en = cfgRegs_17[46]; // @[CGRA.scala 667:42]
  assign gibs_35_io_cfg_addr = cfgRegs_17[45:32]; // @[CGRA.scala 668:44]
  assign gibs_35_io_cfg_data = cfgRegs_17[31:0]; // @[CGRA.scala 669:44]
  assign gibs_35_io_opinNW_0 = pes_23_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_35_io_opinNE_0 = lsus_15_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_35_io_opinSE_0 = lsus_17_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_35_io_opinSW_0 = pes_26_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_35_io_itrackW_0 = gibs_34_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_35_io_itrackN_0 = gibs_31_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_35_io_itrackS_0 = gibs_39_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_36_clock = clock;
  assign gibs_36_reset = reset;
  assign gibs_36_io_cfg_en = cfgRegs_19[46]; // @[CGRA.scala 667:42]
  assign gibs_36_io_cfg_addr = cfgRegs_19[45:32]; // @[CGRA.scala 668:44]
  assign gibs_36_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 669:44]
  assign gibs_36_io_opinNW_0 = lsus_16_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_36_io_opinNE_0 = pes_24_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_36_io_opinSE_0 = pes_27_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_36_io_opinSW_0 = lsus_18_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_36_io_itrackN_0 = gibs_32_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_36_io_itrackE_0 = gibs_37_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_36_io_itrackS_0 = gibs_40_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_37_clock = clock;
  assign gibs_37_reset = reset;
  assign gibs_37_io_cfg_en = cfgRegs_19[46]; // @[CGRA.scala 667:42]
  assign gibs_37_io_cfg_addr = cfgRegs_19[45:32]; // @[CGRA.scala 668:44]
  assign gibs_37_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 669:44]
  assign gibs_37_io_opinNW_0 = pes_24_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_37_io_opinNE_0 = pes_25_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_37_io_opinSE_0 = pes_28_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_37_io_opinSW_0 = pes_27_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_37_io_itrackW_0 = gibs_36_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_37_io_itrackN_0 = gibs_33_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_37_io_itrackE_0 = gibs_38_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_37_io_itrackS_0 = gibs_41_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_38_clock = clock;
  assign gibs_38_reset = reset;
  assign gibs_38_io_cfg_en = cfgRegs_19[46]; // @[CGRA.scala 667:42]
  assign gibs_38_io_cfg_addr = cfgRegs_19[45:32]; // @[CGRA.scala 668:44]
  assign gibs_38_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 669:44]
  assign gibs_38_io_opinNW_0 = pes_25_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_38_io_opinNE_0 = pes_26_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_38_io_opinSE_0 = pes_29_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_38_io_opinSW_0 = pes_28_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_38_io_itrackW_0 = gibs_37_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_38_io_itrackN_0 = gibs_34_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_38_io_itrackE_0 = gibs_39_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_38_io_itrackS_0 = gibs_42_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_39_clock = clock;
  assign gibs_39_reset = reset;
  assign gibs_39_io_cfg_en = cfgRegs_19[46]; // @[CGRA.scala 667:42]
  assign gibs_39_io_cfg_addr = cfgRegs_19[45:32]; // @[CGRA.scala 668:44]
  assign gibs_39_io_cfg_data = cfgRegs_19[31:0]; // @[CGRA.scala 669:44]
  assign gibs_39_io_opinNW_0 = pes_26_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_39_io_opinNE_0 = lsus_17_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_39_io_opinSE_0 = lsus_19_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_39_io_opinSW_0 = pes_29_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_39_io_itrackW_0 = gibs_38_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_39_io_itrackN_0 = gibs_35_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_39_io_itrackS_0 = gibs_43_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_40_clock = clock;
  assign gibs_40_reset = reset;
  assign gibs_40_io_cfg_en = cfgRegs_21[46]; // @[CGRA.scala 667:42]
  assign gibs_40_io_cfg_addr = cfgRegs_21[45:32]; // @[CGRA.scala 668:44]
  assign gibs_40_io_cfg_data = cfgRegs_21[31:0]; // @[CGRA.scala 669:44]
  assign gibs_40_io_opinNW_0 = lsus_18_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_40_io_opinNE_0 = pes_27_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_40_io_opinSE_0 = pes_30_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_40_io_opinSW_0 = lsus_20_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_40_io_itrackN_0 = gibs_36_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_40_io_itrackE_0 = gibs_41_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_40_io_itrackS_0 = gibs_44_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_41_clock = clock;
  assign gibs_41_reset = reset;
  assign gibs_41_io_cfg_en = cfgRegs_21[46]; // @[CGRA.scala 667:42]
  assign gibs_41_io_cfg_addr = cfgRegs_21[45:32]; // @[CGRA.scala 668:44]
  assign gibs_41_io_cfg_data = cfgRegs_21[31:0]; // @[CGRA.scala 669:44]
  assign gibs_41_io_opinNW_0 = pes_27_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_41_io_opinNE_0 = pes_28_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_41_io_opinSE_0 = pes_31_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_41_io_opinSW_0 = pes_30_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_41_io_itrackW_0 = gibs_40_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_41_io_itrackN_0 = gibs_37_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_41_io_itrackE_0 = gibs_42_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_41_io_itrackS_0 = gibs_45_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_42_clock = clock;
  assign gibs_42_reset = reset;
  assign gibs_42_io_cfg_en = cfgRegs_21[46]; // @[CGRA.scala 667:42]
  assign gibs_42_io_cfg_addr = cfgRegs_21[45:32]; // @[CGRA.scala 668:44]
  assign gibs_42_io_cfg_data = cfgRegs_21[31:0]; // @[CGRA.scala 669:44]
  assign gibs_42_io_opinNW_0 = pes_28_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_42_io_opinNE_0 = pes_29_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_42_io_opinSE_0 = pes_32_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_42_io_opinSW_0 = pes_31_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_42_io_itrackW_0 = gibs_41_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_42_io_itrackN_0 = gibs_38_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_42_io_itrackE_0 = gibs_43_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_42_io_itrackS_0 = gibs_46_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_43_clock = clock;
  assign gibs_43_reset = reset;
  assign gibs_43_io_cfg_en = cfgRegs_21[46]; // @[CGRA.scala 667:42]
  assign gibs_43_io_cfg_addr = cfgRegs_21[45:32]; // @[CGRA.scala 668:44]
  assign gibs_43_io_cfg_data = cfgRegs_21[31:0]; // @[CGRA.scala 669:44]
  assign gibs_43_io_opinNW_0 = pes_29_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_43_io_opinNE_0 = lsus_19_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_43_io_opinSE_0 = lsus_21_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_43_io_opinSW_0 = pes_32_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_43_io_itrackW_0 = gibs_42_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_43_io_itrackN_0 = gibs_39_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_43_io_itrackS_0 = gibs_47_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_44_clock = clock;
  assign gibs_44_reset = reset;
  assign gibs_44_io_cfg_en = cfgRegs_23[46]; // @[CGRA.scala 667:42]
  assign gibs_44_io_cfg_addr = cfgRegs_23[45:32]; // @[CGRA.scala 668:44]
  assign gibs_44_io_cfg_data = cfgRegs_23[31:0]; // @[CGRA.scala 669:44]
  assign gibs_44_io_opinNW_0 = lsus_20_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_44_io_opinNE_0 = pes_30_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_44_io_opinSE_0 = pes_33_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_44_io_opinSW_0 = lsus_22_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_44_io_itrackN_0 = gibs_40_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_44_io_itrackE_0 = gibs_45_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_44_io_itrackS_0 = gibs_48_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_45_clock = clock;
  assign gibs_45_reset = reset;
  assign gibs_45_io_cfg_en = cfgRegs_23[46]; // @[CGRA.scala 667:42]
  assign gibs_45_io_cfg_addr = cfgRegs_23[45:32]; // @[CGRA.scala 668:44]
  assign gibs_45_io_cfg_data = cfgRegs_23[31:0]; // @[CGRA.scala 669:44]
  assign gibs_45_io_opinNW_0 = pes_30_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_45_io_opinNE_0 = pes_31_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_45_io_opinSE_0 = pes_34_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_45_io_opinSW_0 = pes_33_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_45_io_itrackW_0 = gibs_44_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_45_io_itrackN_0 = gibs_41_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_45_io_itrackE_0 = gibs_46_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_45_io_itrackS_0 = gibs_49_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_46_clock = clock;
  assign gibs_46_reset = reset;
  assign gibs_46_io_cfg_en = cfgRegs_23[46]; // @[CGRA.scala 667:42]
  assign gibs_46_io_cfg_addr = cfgRegs_23[45:32]; // @[CGRA.scala 668:44]
  assign gibs_46_io_cfg_data = cfgRegs_23[31:0]; // @[CGRA.scala 669:44]
  assign gibs_46_io_opinNW_0 = pes_31_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_46_io_opinNE_0 = pes_32_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_46_io_opinSE_0 = pes_35_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_46_io_opinSW_0 = pes_34_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_46_io_itrackW_0 = gibs_45_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_46_io_itrackN_0 = gibs_42_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_46_io_itrackE_0 = gibs_47_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_46_io_itrackS_0 = gibs_50_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_47_clock = clock;
  assign gibs_47_reset = reset;
  assign gibs_47_io_cfg_en = cfgRegs_23[46]; // @[CGRA.scala 667:42]
  assign gibs_47_io_cfg_addr = cfgRegs_23[45:32]; // @[CGRA.scala 668:44]
  assign gibs_47_io_cfg_data = cfgRegs_23[31:0]; // @[CGRA.scala 669:44]
  assign gibs_47_io_opinNW_0 = pes_32_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_47_io_opinNE_0 = lsus_21_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_47_io_opinSE_0 = lsus_23_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_47_io_opinSW_0 = pes_35_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_47_io_itrackW_0 = gibs_46_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_47_io_itrackN_0 = gibs_43_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_47_io_itrackS_0 = gibs_51_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_48_clock = clock;
  assign gibs_48_reset = reset;
  assign gibs_48_io_cfg_en = cfgRegs_25[46]; // @[CGRA.scala 667:42]
  assign gibs_48_io_cfg_addr = cfgRegs_25[45:32]; // @[CGRA.scala 668:44]
  assign gibs_48_io_cfg_data = cfgRegs_25[31:0]; // @[CGRA.scala 669:44]
  assign gibs_48_io_opinNW_0 = lsus_22_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_48_io_opinNE_0 = pes_33_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_48_io_opinSE_0 = pes_36_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_48_io_opinSW_0 = lsus_24_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_48_io_itrackN_0 = gibs_44_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_48_io_itrackE_0 = gibs_49_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_48_io_itrackS_0 = gibs_52_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_49_clock = clock;
  assign gibs_49_reset = reset;
  assign gibs_49_io_cfg_en = cfgRegs_25[46]; // @[CGRA.scala 667:42]
  assign gibs_49_io_cfg_addr = cfgRegs_25[45:32]; // @[CGRA.scala 668:44]
  assign gibs_49_io_cfg_data = cfgRegs_25[31:0]; // @[CGRA.scala 669:44]
  assign gibs_49_io_opinNW_0 = pes_33_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_49_io_opinNE_0 = pes_34_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_49_io_opinSE_0 = pes_37_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_49_io_opinSW_0 = pes_36_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_49_io_itrackW_0 = gibs_48_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_49_io_itrackN_0 = gibs_45_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_49_io_itrackE_0 = gibs_50_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_49_io_itrackS_0 = gibs_53_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_50_clock = clock;
  assign gibs_50_reset = reset;
  assign gibs_50_io_cfg_en = cfgRegs_25[46]; // @[CGRA.scala 667:42]
  assign gibs_50_io_cfg_addr = cfgRegs_25[45:32]; // @[CGRA.scala 668:44]
  assign gibs_50_io_cfg_data = cfgRegs_25[31:0]; // @[CGRA.scala 669:44]
  assign gibs_50_io_opinNW_0 = pes_34_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_50_io_opinNE_0 = pes_35_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_50_io_opinSE_0 = pes_38_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_50_io_opinSW_0 = pes_37_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_50_io_itrackW_0 = gibs_49_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_50_io_itrackN_0 = gibs_46_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_50_io_itrackE_0 = gibs_51_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_50_io_itrackS_0 = gibs_54_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_51_clock = clock;
  assign gibs_51_reset = reset;
  assign gibs_51_io_cfg_en = cfgRegs_25[46]; // @[CGRA.scala 667:42]
  assign gibs_51_io_cfg_addr = cfgRegs_25[45:32]; // @[CGRA.scala 668:44]
  assign gibs_51_io_cfg_data = cfgRegs_25[31:0]; // @[CGRA.scala 669:44]
  assign gibs_51_io_opinNW_0 = pes_35_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_51_io_opinNE_0 = lsus_23_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_51_io_opinSE_0 = lsus_25_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_51_io_opinSW_0 = pes_38_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_51_io_itrackW_0 = gibs_50_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_51_io_itrackN_0 = gibs_47_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_51_io_itrackS_0 = gibs_55_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_52_clock = clock;
  assign gibs_52_reset = reset;
  assign gibs_52_io_cfg_en = cfgRegs_27[46]; // @[CGRA.scala 667:42]
  assign gibs_52_io_cfg_addr = cfgRegs_27[45:32]; // @[CGRA.scala 668:44]
  assign gibs_52_io_cfg_data = cfgRegs_27[31:0]; // @[CGRA.scala 669:44]
  assign gibs_52_io_opinNW_0 = lsus_24_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_52_io_opinNE_0 = pes_36_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_52_io_opinSE_0 = pes_39_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_52_io_opinSW_0 = lsus_26_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_52_io_itrackN_0 = gibs_48_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_52_io_itrackE_0 = gibs_53_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_52_io_itrackS_0 = gibs_56_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_53_clock = clock;
  assign gibs_53_reset = reset;
  assign gibs_53_io_cfg_en = cfgRegs_27[46]; // @[CGRA.scala 667:42]
  assign gibs_53_io_cfg_addr = cfgRegs_27[45:32]; // @[CGRA.scala 668:44]
  assign gibs_53_io_cfg_data = cfgRegs_27[31:0]; // @[CGRA.scala 669:44]
  assign gibs_53_io_opinNW_0 = pes_36_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_53_io_opinNE_0 = pes_37_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_53_io_opinSE_0 = pes_40_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_53_io_opinSW_0 = pes_39_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_53_io_itrackW_0 = gibs_52_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_53_io_itrackN_0 = gibs_49_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_53_io_itrackE_0 = gibs_54_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_53_io_itrackS_0 = gibs_57_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_54_clock = clock;
  assign gibs_54_reset = reset;
  assign gibs_54_io_cfg_en = cfgRegs_27[46]; // @[CGRA.scala 667:42]
  assign gibs_54_io_cfg_addr = cfgRegs_27[45:32]; // @[CGRA.scala 668:44]
  assign gibs_54_io_cfg_data = cfgRegs_27[31:0]; // @[CGRA.scala 669:44]
  assign gibs_54_io_opinNW_0 = pes_37_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_54_io_opinNE_0 = pes_38_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_54_io_opinSE_0 = pes_41_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_54_io_opinSW_0 = pes_40_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_54_io_itrackW_0 = gibs_53_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_54_io_itrackN_0 = gibs_50_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_54_io_itrackE_0 = gibs_55_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_54_io_itrackS_0 = gibs_58_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_55_clock = clock;
  assign gibs_55_reset = reset;
  assign gibs_55_io_cfg_en = cfgRegs_27[46]; // @[CGRA.scala 667:42]
  assign gibs_55_io_cfg_addr = cfgRegs_27[45:32]; // @[CGRA.scala 668:44]
  assign gibs_55_io_cfg_data = cfgRegs_27[31:0]; // @[CGRA.scala 669:44]
  assign gibs_55_io_opinNW_0 = pes_38_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_55_io_opinNE_0 = lsus_25_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_55_io_opinSE_0 = lsus_27_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_55_io_opinSW_0 = pes_41_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_55_io_itrackW_0 = gibs_54_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_55_io_itrackN_0 = gibs_51_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_55_io_itrackS_0 = gibs_59_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_56_clock = clock;
  assign gibs_56_reset = reset;
  assign gibs_56_io_cfg_en = cfgRegs_29[46]; // @[CGRA.scala 667:42]
  assign gibs_56_io_cfg_addr = cfgRegs_29[45:32]; // @[CGRA.scala 668:44]
  assign gibs_56_io_cfg_data = cfgRegs_29[31:0]; // @[CGRA.scala 669:44]
  assign gibs_56_io_opinNW_0 = lsus_26_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_56_io_opinNE_0 = pes_39_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_56_io_opinSE_0 = pes_42_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_56_io_opinSW_0 = lsus_28_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_56_io_itrackN_0 = gibs_52_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_56_io_itrackE_0 = gibs_57_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_56_io_itrackS_0 = gibs_60_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_57_clock = clock;
  assign gibs_57_reset = reset;
  assign gibs_57_io_cfg_en = cfgRegs_29[46]; // @[CGRA.scala 667:42]
  assign gibs_57_io_cfg_addr = cfgRegs_29[45:32]; // @[CGRA.scala 668:44]
  assign gibs_57_io_cfg_data = cfgRegs_29[31:0]; // @[CGRA.scala 669:44]
  assign gibs_57_io_opinNW_0 = pes_39_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_57_io_opinNE_0 = pes_40_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_57_io_opinSE_0 = pes_43_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_57_io_opinSW_0 = pes_42_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_57_io_itrackW_0 = gibs_56_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_57_io_itrackN_0 = gibs_53_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_57_io_itrackE_0 = gibs_58_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_57_io_itrackS_0 = gibs_61_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_58_clock = clock;
  assign gibs_58_reset = reset;
  assign gibs_58_io_cfg_en = cfgRegs_29[46]; // @[CGRA.scala 667:42]
  assign gibs_58_io_cfg_addr = cfgRegs_29[45:32]; // @[CGRA.scala 668:44]
  assign gibs_58_io_cfg_data = cfgRegs_29[31:0]; // @[CGRA.scala 669:44]
  assign gibs_58_io_opinNW_0 = pes_40_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_58_io_opinNE_0 = pes_41_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_58_io_opinSE_0 = pes_44_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_58_io_opinSW_0 = pes_43_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_58_io_itrackW_0 = gibs_57_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_58_io_itrackN_0 = gibs_54_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_58_io_itrackE_0 = gibs_59_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_58_io_itrackS_0 = gibs_62_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_59_clock = clock;
  assign gibs_59_reset = reset;
  assign gibs_59_io_cfg_en = cfgRegs_29[46]; // @[CGRA.scala 667:42]
  assign gibs_59_io_cfg_addr = cfgRegs_29[45:32]; // @[CGRA.scala 668:44]
  assign gibs_59_io_cfg_data = cfgRegs_29[31:0]; // @[CGRA.scala 669:44]
  assign gibs_59_io_opinNW_0 = pes_41_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_59_io_opinNE_0 = lsus_27_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_59_io_opinSE_0 = lsus_29_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_59_io_opinSW_0 = pes_44_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_59_io_itrackW_0 = gibs_58_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_59_io_itrackN_0 = gibs_55_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_59_io_itrackS_0 = gibs_63_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_60_clock = clock;
  assign gibs_60_reset = reset;
  assign gibs_60_io_cfg_en = cfgRegs_31[46]; // @[CGRA.scala 667:42]
  assign gibs_60_io_cfg_addr = cfgRegs_31[45:32]; // @[CGRA.scala 668:44]
  assign gibs_60_io_cfg_data = cfgRegs_31[31:0]; // @[CGRA.scala 669:44]
  assign gibs_60_io_opinNW_0 = lsus_28_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_60_io_opinNE_0 = pes_42_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_60_io_opinSE_0 = pes_45_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_60_io_opinSW_0 = lsus_30_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_60_io_itrackN_0 = gibs_56_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_60_io_itrackE_0 = gibs_61_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_60_io_itrackS_0 = gibs_64_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_61_clock = clock;
  assign gibs_61_reset = reset;
  assign gibs_61_io_cfg_en = cfgRegs_31[46]; // @[CGRA.scala 667:42]
  assign gibs_61_io_cfg_addr = cfgRegs_31[45:32]; // @[CGRA.scala 668:44]
  assign gibs_61_io_cfg_data = cfgRegs_31[31:0]; // @[CGRA.scala 669:44]
  assign gibs_61_io_opinNW_0 = pes_42_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_61_io_opinNE_0 = pes_43_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_61_io_opinSE_0 = pes_46_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_61_io_opinSW_0 = pes_45_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_61_io_itrackW_0 = gibs_60_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_61_io_itrackN_0 = gibs_57_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_61_io_itrackE_0 = gibs_62_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_61_io_itrackS_0 = gibs_65_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_62_clock = clock;
  assign gibs_62_reset = reset;
  assign gibs_62_io_cfg_en = cfgRegs_31[46]; // @[CGRA.scala 667:42]
  assign gibs_62_io_cfg_addr = cfgRegs_31[45:32]; // @[CGRA.scala 668:44]
  assign gibs_62_io_cfg_data = cfgRegs_31[31:0]; // @[CGRA.scala 669:44]
  assign gibs_62_io_opinNW_0 = pes_43_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_62_io_opinNE_0 = pes_44_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_62_io_opinSE_0 = pes_47_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_62_io_opinSW_0 = pes_46_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_62_io_itrackW_0 = gibs_61_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_62_io_itrackN_0 = gibs_58_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_62_io_itrackE_0 = gibs_63_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_62_io_itrackS_0 = gibs_66_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_63_clock = clock;
  assign gibs_63_reset = reset;
  assign gibs_63_io_cfg_en = cfgRegs_31[46]; // @[CGRA.scala 667:42]
  assign gibs_63_io_cfg_addr = cfgRegs_31[45:32]; // @[CGRA.scala 668:44]
  assign gibs_63_io_cfg_data = cfgRegs_31[31:0]; // @[CGRA.scala 669:44]
  assign gibs_63_io_opinNW_0 = pes_44_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_63_io_opinNE_0 = lsus_29_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_63_io_opinSE_0 = lsus_31_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_63_io_opinSW_0 = pes_47_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_63_io_itrackW_0 = gibs_62_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_63_io_itrackN_0 = gibs_59_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_63_io_itrackS_0 = gibs_67_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_64_clock = clock;
  assign gibs_64_reset = reset;
  assign gibs_64_io_cfg_en = cfgRegs_33[46]; // @[CGRA.scala 667:42]
  assign gibs_64_io_cfg_addr = cfgRegs_33[45:32]; // @[CGRA.scala 668:44]
  assign gibs_64_io_cfg_data = cfgRegs_33[31:0]; // @[CGRA.scala 669:44]
  assign gibs_64_io_opinNW_0 = lsus_30_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_64_io_opinNE_0 = pes_45_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_64_io_opinSE_0 = pes_48_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_64_io_opinSW_0 = lsus_32_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_64_io_itrackN_0 = gibs_60_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_64_io_itrackE_0 = gibs_65_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_64_io_itrackS_0 = gibs_68_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_65_clock = clock;
  assign gibs_65_reset = reset;
  assign gibs_65_io_cfg_en = cfgRegs_33[46]; // @[CGRA.scala 667:42]
  assign gibs_65_io_cfg_addr = cfgRegs_33[45:32]; // @[CGRA.scala 668:44]
  assign gibs_65_io_cfg_data = cfgRegs_33[31:0]; // @[CGRA.scala 669:44]
  assign gibs_65_io_opinNW_0 = pes_45_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_65_io_opinNE_0 = pes_46_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_65_io_opinSE_0 = pes_49_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_65_io_opinSW_0 = pes_48_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_65_io_itrackW_0 = gibs_64_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_65_io_itrackN_0 = gibs_61_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_65_io_itrackE_0 = gibs_66_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_65_io_itrackS_0 = gibs_69_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_66_clock = clock;
  assign gibs_66_reset = reset;
  assign gibs_66_io_cfg_en = cfgRegs_33[46]; // @[CGRA.scala 667:42]
  assign gibs_66_io_cfg_addr = cfgRegs_33[45:32]; // @[CGRA.scala 668:44]
  assign gibs_66_io_cfg_data = cfgRegs_33[31:0]; // @[CGRA.scala 669:44]
  assign gibs_66_io_opinNW_0 = pes_46_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_66_io_opinNE_0 = pes_47_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_66_io_opinSE_0 = pes_50_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_66_io_opinSW_0 = pes_49_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_66_io_itrackW_0 = gibs_65_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_66_io_itrackN_0 = gibs_62_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_66_io_itrackE_0 = gibs_67_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_66_io_itrackS_0 = gibs_70_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_67_clock = clock;
  assign gibs_67_reset = reset;
  assign gibs_67_io_cfg_en = cfgRegs_33[46]; // @[CGRA.scala 667:42]
  assign gibs_67_io_cfg_addr = cfgRegs_33[45:32]; // @[CGRA.scala 668:44]
  assign gibs_67_io_cfg_data = cfgRegs_33[31:0]; // @[CGRA.scala 669:44]
  assign gibs_67_io_opinNW_0 = pes_47_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_67_io_opinNE_0 = lsus_31_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_67_io_opinSE_0 = lsus_33_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_67_io_opinSW_0 = pes_50_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_67_io_itrackW_0 = gibs_66_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_67_io_itrackN_0 = gibs_63_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_67_io_itrackS_0 = gibs_71_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_68_clock = clock;
  assign gibs_68_reset = reset;
  assign gibs_68_io_cfg_en = cfgRegs_35[46]; // @[CGRA.scala 667:42]
  assign gibs_68_io_cfg_addr = cfgRegs_35[45:32]; // @[CGRA.scala 668:44]
  assign gibs_68_io_cfg_data = cfgRegs_35[31:0]; // @[CGRA.scala 669:44]
  assign gibs_68_io_opinNW_0 = lsus_32_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_68_io_opinNE_0 = pes_48_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_68_io_opinSE_0 = pes_51_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_68_io_opinSW_0 = lsus_34_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_68_io_itrackN_0 = gibs_64_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_68_io_itrackE_0 = gibs_69_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_68_io_itrackS_0 = gibs_72_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_69_clock = clock;
  assign gibs_69_reset = reset;
  assign gibs_69_io_cfg_en = cfgRegs_35[46]; // @[CGRA.scala 667:42]
  assign gibs_69_io_cfg_addr = cfgRegs_35[45:32]; // @[CGRA.scala 668:44]
  assign gibs_69_io_cfg_data = cfgRegs_35[31:0]; // @[CGRA.scala 669:44]
  assign gibs_69_io_opinNW_0 = pes_48_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_69_io_opinNE_0 = pes_49_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_69_io_opinSE_0 = pes_52_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_69_io_opinSW_0 = pes_51_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_69_io_itrackW_0 = gibs_68_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_69_io_itrackN_0 = gibs_65_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_69_io_itrackE_0 = gibs_70_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_69_io_itrackS_0 = gibs_73_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_70_clock = clock;
  assign gibs_70_reset = reset;
  assign gibs_70_io_cfg_en = cfgRegs_35[46]; // @[CGRA.scala 667:42]
  assign gibs_70_io_cfg_addr = cfgRegs_35[45:32]; // @[CGRA.scala 668:44]
  assign gibs_70_io_cfg_data = cfgRegs_35[31:0]; // @[CGRA.scala 669:44]
  assign gibs_70_io_opinNW_0 = pes_49_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_70_io_opinNE_0 = pes_50_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_70_io_opinSE_0 = pes_53_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_70_io_opinSW_0 = pes_52_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_70_io_itrackW_0 = gibs_69_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_70_io_itrackN_0 = gibs_66_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_70_io_itrackE_0 = gibs_71_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_70_io_itrackS_0 = gibs_74_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_71_clock = clock;
  assign gibs_71_reset = reset;
  assign gibs_71_io_cfg_en = cfgRegs_35[46]; // @[CGRA.scala 667:42]
  assign gibs_71_io_cfg_addr = cfgRegs_35[45:32]; // @[CGRA.scala 668:44]
  assign gibs_71_io_cfg_data = cfgRegs_35[31:0]; // @[CGRA.scala 669:44]
  assign gibs_71_io_opinNW_0 = pes_50_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_71_io_opinNE_0 = lsus_33_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_71_io_opinSE_0 = lsus_35_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_71_io_opinSW_0 = pes_53_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_71_io_itrackW_0 = gibs_70_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_71_io_itrackN_0 = gibs_67_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_71_io_itrackS_0 = gibs_75_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_72_clock = clock;
  assign gibs_72_reset = reset;
  assign gibs_72_io_cfg_en = cfgRegs_37[46]; // @[CGRA.scala 667:42]
  assign gibs_72_io_cfg_addr = cfgRegs_37[45:32]; // @[CGRA.scala 668:44]
  assign gibs_72_io_cfg_data = cfgRegs_37[31:0]; // @[CGRA.scala 669:44]
  assign gibs_72_io_opinNW_0 = lsus_34_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_72_io_opinNE_0 = pes_51_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_72_io_opinSE_0 = pes_54_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_72_io_opinSW_0 = lsus_36_io_out_0; // @[CGRA.scala 609:39]
  assign gibs_72_io_itrackN_0 = gibs_68_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_72_io_itrackE_0 = gibs_73_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_72_io_itrackS_0 = gibs_76_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_73_clock = clock;
  assign gibs_73_reset = reset;
  assign gibs_73_io_cfg_en = cfgRegs_37[46]; // @[CGRA.scala 667:42]
  assign gibs_73_io_cfg_addr = cfgRegs_37[45:32]; // @[CGRA.scala 668:44]
  assign gibs_73_io_cfg_data = cfgRegs_37[31:0]; // @[CGRA.scala 669:44]
  assign gibs_73_io_opinNW_0 = pes_51_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_73_io_opinNE_0 = pes_52_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_73_io_opinSE_0 = pes_55_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_73_io_opinSW_0 = pes_54_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_73_io_itrackW_0 = gibs_72_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_73_io_itrackN_0 = gibs_69_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_73_io_itrackE_0 = gibs_74_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_73_io_itrackS_0 = gibs_77_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_74_clock = clock;
  assign gibs_74_reset = reset;
  assign gibs_74_io_cfg_en = cfgRegs_37[46]; // @[CGRA.scala 667:42]
  assign gibs_74_io_cfg_addr = cfgRegs_37[45:32]; // @[CGRA.scala 668:44]
  assign gibs_74_io_cfg_data = cfgRegs_37[31:0]; // @[CGRA.scala 669:44]
  assign gibs_74_io_opinNW_0 = pes_52_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_74_io_opinNE_0 = pes_53_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_74_io_opinSE_0 = pes_56_io_out_0; // @[CGRA.scala 497:41]
  assign gibs_74_io_opinSW_0 = pes_55_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_74_io_itrackW_0 = gibs_73_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_74_io_itrackN_0 = gibs_70_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_74_io_itrackE_0 = gibs_75_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_74_io_itrackS_0 = gibs_78_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_75_clock = clock;
  assign gibs_75_reset = reset;
  assign gibs_75_io_cfg_en = cfgRegs_37[46]; // @[CGRA.scala 667:42]
  assign gibs_75_io_cfg_addr = cfgRegs_37[45:32]; // @[CGRA.scala 668:44]
  assign gibs_75_io_cfg_data = cfgRegs_37[31:0]; // @[CGRA.scala 669:44]
  assign gibs_75_io_opinNW_0 = pes_53_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_75_io_opinNE_0 = lsus_35_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_75_io_opinSE_0 = lsus_37_io_out_0; // @[CGRA.scala 629:46]
  assign gibs_75_io_opinSW_0 = pes_56_io_out_0; // @[CGRA.scala 498:43]
  assign gibs_75_io_itrackW_0 = gibs_74_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_75_io_itrackN_0 = gibs_71_io_otrackS_0; // @[CGRA.scala 538:16]
  assign gibs_75_io_itrackS_0 = gibs_79_io_otrackN_0; // @[CGRA.scala 544:16]
  assign gibs_76_clock = clock;
  assign gibs_76_reset = reset;
  assign gibs_76_io_cfg_en = cfgRegs_39[46]; // @[CGRA.scala 667:42]
  assign gibs_76_io_cfg_addr = cfgRegs_39[45:32]; // @[CGRA.scala 668:44]
  assign gibs_76_io_cfg_data = cfgRegs_39[31:0]; // @[CGRA.scala 669:44]
  assign gibs_76_io_opinNW_0 = lsus_36_io_out_0; // @[CGRA.scala 610:43]
  assign gibs_76_io_opinNE_0 = pes_54_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_76_io_opinSE_0 = ibs_3_io_out_0; // @[CGRA.scala 428:35]
  assign gibs_76_io_itrackN_0 = gibs_72_io_otrackS_0; // @[CGRA.scala 530:16]
  assign gibs_76_io_itrackE_0 = gibs_77_io_otrackW_0; // @[CGRA.scala 554:16]
  assign gibs_77_clock = clock;
  assign gibs_77_reset = reset;
  assign gibs_77_io_cfg_en = cfgRegs_39[46]; // @[CGRA.scala 667:42]
  assign gibs_77_io_cfg_addr = cfgRegs_39[45:32]; // @[CGRA.scala 668:44]
  assign gibs_77_io_cfg_data = cfgRegs_39[31:0]; // @[CGRA.scala 669:44]
  assign gibs_77_io_opinNW_0 = pes_54_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_77_io_opinNE_0 = pes_55_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_77_io_opinSE_0 = ibs_4_io_out_0; // @[CGRA.scala 428:35]
  assign gibs_77_io_opinSW_0 = ibs_3_io_out_0; // @[CGRA.scala 429:37]
  assign gibs_77_io_itrackW_0 = gibs_76_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_77_io_itrackN_0 = gibs_73_io_otrackS_0; // @[CGRA.scala 530:16]
  assign gibs_77_io_itrackE_0 = gibs_78_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_78_clock = clock;
  assign gibs_78_reset = reset;
  assign gibs_78_io_cfg_en = cfgRegs_39[46]; // @[CGRA.scala 667:42]
  assign gibs_78_io_cfg_addr = cfgRegs_39[45:32]; // @[CGRA.scala 668:44]
  assign gibs_78_io_cfg_data = cfgRegs_39[31:0]; // @[CGRA.scala 669:44]
  assign gibs_78_io_opinNW_0 = pes_55_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_78_io_opinNE_0 = pes_56_io_out_0; // @[CGRA.scala 499:45]
  assign gibs_78_io_opinSE_0 = ibs_5_io_out_0; // @[CGRA.scala 428:35]
  assign gibs_78_io_opinSW_0 = ibs_4_io_out_0; // @[CGRA.scala 429:37]
  assign gibs_78_io_itrackW_0 = gibs_77_io_otrackE_0; // @[CGRA.scala 571:16]
  assign gibs_78_io_itrackN_0 = gibs_74_io_otrackS_0; // @[CGRA.scala 530:16]
  assign gibs_78_io_itrackE_0 = gibs_79_io_otrackW_0; // @[CGRA.scala 577:16]
  assign gibs_79_clock = clock;
  assign gibs_79_reset = reset;
  assign gibs_79_io_cfg_en = cfgRegs_39[46]; // @[CGRA.scala 667:42]
  assign gibs_79_io_cfg_addr = cfgRegs_39[45:32]; // @[CGRA.scala 668:44]
  assign gibs_79_io_cfg_data = cfgRegs_39[31:0]; // @[CGRA.scala 669:44]
  assign gibs_79_io_opinNW_0 = pes_56_io_out_0; // @[CGRA.scala 500:47]
  assign gibs_79_io_opinNE_0 = lsus_37_io_out_0; // @[CGRA.scala 630:50]
  assign gibs_79_io_opinSW_0 = ibs_5_io_out_0; // @[CGRA.scala 429:37]
  assign gibs_79_io_itrackW_0 = gibs_78_io_otrackE_0; // @[CGRA.scala 563:16]
  assign gibs_79_io_itrackN_0 = gibs_75_io_otrackS_0; // @[CGRA.scala 530:16]
  assign lsus_0_clock = clock;
  assign lsus_0_reset = reset;
  assign lsus_0_io_cfg_en = cfgRegs_2[46]; // @[CGRA.scala 678:35]
  assign lsus_0_io_cfg_addr = cfgRegs_2[45:32]; // @[CGRA.scala 679:37]
  assign lsus_0_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 680:37]
  assign lsus_0_io_hostInterface_read_addr = io_hostInterface_0_read_addr; // @[CGRA.scala 595:36]
  assign lsus_0_io_hostInterface_read_data_ready = io_hostInterface_0_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_0_io_hostInterface_write_addr = io_hostInterface_0_write_addr; // @[CGRA.scala 595:36]
  assign lsus_0_io_hostInterface_write_data_valid = io_hostInterface_0_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_0_io_hostInterface_write_data_bits = io_hostInterface_0_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_0_io_hostInterface_cycle = io_hostInterface_0_cycle; // @[CGRA.scala 595:36]
  assign lsus_0_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_0_io_in_0 = gibs_0_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_0_io_in_1 = gibs_4_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_1_clock = clock;
  assign lsus_1_reset = reset;
  assign lsus_1_io_cfg_en = cfgRegs_2[46]; // @[CGRA.scala 678:35]
  assign lsus_1_io_cfg_addr = cfgRegs_2[45:32]; // @[CGRA.scala 679:37]
  assign lsus_1_io_cfg_data = cfgRegs_2[31:0]; // @[CGRA.scala 680:37]
  assign lsus_1_io_hostInterface_read_addr = io_hostInterface_1_read_addr; // @[CGRA.scala 595:36]
  assign lsus_1_io_hostInterface_read_data_ready = io_hostInterface_1_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_1_io_hostInterface_write_addr = io_hostInterface_1_write_addr; // @[CGRA.scala 595:36]
  assign lsus_1_io_hostInterface_write_data_valid = io_hostInterface_1_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_1_io_hostInterface_write_data_bits = io_hostInterface_1_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_1_io_hostInterface_cycle = io_hostInterface_1_cycle; // @[CGRA.scala 595:36]
  assign lsus_1_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_1_io_in_0 = gibs_3_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_1_io_in_1 = gibs_7_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_2_clock = clock;
  assign lsus_2_reset = reset;
  assign lsus_2_io_cfg_en = cfgRegs_4[46]; // @[CGRA.scala 678:35]
  assign lsus_2_io_cfg_addr = cfgRegs_4[45:32]; // @[CGRA.scala 679:37]
  assign lsus_2_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 680:37]
  assign lsus_2_io_hostInterface_read_addr = io_hostInterface_2_read_addr; // @[CGRA.scala 595:36]
  assign lsus_2_io_hostInterface_read_data_ready = io_hostInterface_2_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_2_io_hostInterface_write_addr = io_hostInterface_2_write_addr; // @[CGRA.scala 595:36]
  assign lsus_2_io_hostInterface_write_data_valid = io_hostInterface_2_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_2_io_hostInterface_write_data_bits = io_hostInterface_2_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_2_io_hostInterface_cycle = io_hostInterface_2_cycle; // @[CGRA.scala 595:36]
  assign lsus_2_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_2_io_in_0 = gibs_4_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_2_io_in_1 = gibs_8_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_3_clock = clock;
  assign lsus_3_reset = reset;
  assign lsus_3_io_cfg_en = cfgRegs_4[46]; // @[CGRA.scala 678:35]
  assign lsus_3_io_cfg_addr = cfgRegs_4[45:32]; // @[CGRA.scala 679:37]
  assign lsus_3_io_cfg_data = cfgRegs_4[31:0]; // @[CGRA.scala 680:37]
  assign lsus_3_io_hostInterface_read_addr = io_hostInterface_3_read_addr; // @[CGRA.scala 595:36]
  assign lsus_3_io_hostInterface_read_data_ready = io_hostInterface_3_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_3_io_hostInterface_write_addr = io_hostInterface_3_write_addr; // @[CGRA.scala 595:36]
  assign lsus_3_io_hostInterface_write_data_valid = io_hostInterface_3_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_3_io_hostInterface_write_data_bits = io_hostInterface_3_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_3_io_hostInterface_cycle = io_hostInterface_3_cycle; // @[CGRA.scala 595:36]
  assign lsus_3_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_3_io_in_0 = gibs_7_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_3_io_in_1 = gibs_11_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_4_clock = clock;
  assign lsus_4_reset = reset;
  assign lsus_4_io_cfg_en = cfgRegs_6[46]; // @[CGRA.scala 678:35]
  assign lsus_4_io_cfg_addr = cfgRegs_6[45:32]; // @[CGRA.scala 679:37]
  assign lsus_4_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 680:37]
  assign lsus_4_io_hostInterface_read_addr = io_hostInterface_4_read_addr; // @[CGRA.scala 595:36]
  assign lsus_4_io_hostInterface_read_data_ready = io_hostInterface_4_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_4_io_hostInterface_write_addr = io_hostInterface_4_write_addr; // @[CGRA.scala 595:36]
  assign lsus_4_io_hostInterface_write_data_valid = io_hostInterface_4_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_4_io_hostInterface_write_data_bits = io_hostInterface_4_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_4_io_hostInterface_cycle = io_hostInterface_4_cycle; // @[CGRA.scala 595:36]
  assign lsus_4_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_4_io_in_0 = gibs_8_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_4_io_in_1 = gibs_12_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_5_clock = clock;
  assign lsus_5_reset = reset;
  assign lsus_5_io_cfg_en = cfgRegs_6[46]; // @[CGRA.scala 678:35]
  assign lsus_5_io_cfg_addr = cfgRegs_6[45:32]; // @[CGRA.scala 679:37]
  assign lsus_5_io_cfg_data = cfgRegs_6[31:0]; // @[CGRA.scala 680:37]
  assign lsus_5_io_hostInterface_read_addr = io_hostInterface_5_read_addr; // @[CGRA.scala 595:36]
  assign lsus_5_io_hostInterface_read_data_ready = io_hostInterface_5_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_5_io_hostInterface_write_addr = io_hostInterface_5_write_addr; // @[CGRA.scala 595:36]
  assign lsus_5_io_hostInterface_write_data_valid = io_hostInterface_5_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_5_io_hostInterface_write_data_bits = io_hostInterface_5_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_5_io_hostInterface_cycle = io_hostInterface_5_cycle; // @[CGRA.scala 595:36]
  assign lsus_5_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_5_io_in_0 = gibs_11_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_5_io_in_1 = gibs_15_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_6_clock = clock;
  assign lsus_6_reset = reset;
  assign lsus_6_io_cfg_en = cfgRegs_8[46]; // @[CGRA.scala 678:35]
  assign lsus_6_io_cfg_addr = cfgRegs_8[45:32]; // @[CGRA.scala 679:37]
  assign lsus_6_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 680:37]
  assign lsus_6_io_hostInterface_read_addr = io_hostInterface_6_read_addr; // @[CGRA.scala 595:36]
  assign lsus_6_io_hostInterface_read_data_ready = io_hostInterface_6_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_6_io_hostInterface_write_addr = io_hostInterface_6_write_addr; // @[CGRA.scala 595:36]
  assign lsus_6_io_hostInterface_write_data_valid = io_hostInterface_6_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_6_io_hostInterface_write_data_bits = io_hostInterface_6_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_6_io_hostInterface_cycle = io_hostInterface_6_cycle; // @[CGRA.scala 595:36]
  assign lsus_6_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_6_io_in_0 = gibs_12_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_6_io_in_1 = gibs_16_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_7_clock = clock;
  assign lsus_7_reset = reset;
  assign lsus_7_io_cfg_en = cfgRegs_8[46]; // @[CGRA.scala 678:35]
  assign lsus_7_io_cfg_addr = cfgRegs_8[45:32]; // @[CGRA.scala 679:37]
  assign lsus_7_io_cfg_data = cfgRegs_8[31:0]; // @[CGRA.scala 680:37]
  assign lsus_7_io_hostInterface_read_addr = io_hostInterface_7_read_addr; // @[CGRA.scala 595:36]
  assign lsus_7_io_hostInterface_read_data_ready = io_hostInterface_7_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_7_io_hostInterface_write_addr = io_hostInterface_7_write_addr; // @[CGRA.scala 595:36]
  assign lsus_7_io_hostInterface_write_data_valid = io_hostInterface_7_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_7_io_hostInterface_write_data_bits = io_hostInterface_7_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_7_io_hostInterface_cycle = io_hostInterface_7_cycle; // @[CGRA.scala 595:36]
  assign lsus_7_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_7_io_in_0 = gibs_15_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_7_io_in_1 = gibs_19_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_8_clock = clock;
  assign lsus_8_reset = reset;
  assign lsus_8_io_cfg_en = cfgRegs_10[46]; // @[CGRA.scala 678:35]
  assign lsus_8_io_cfg_addr = cfgRegs_10[45:32]; // @[CGRA.scala 679:37]
  assign lsus_8_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 680:37]
  assign lsus_8_io_hostInterface_read_addr = io_hostInterface_8_read_addr; // @[CGRA.scala 595:36]
  assign lsus_8_io_hostInterface_read_data_ready = io_hostInterface_8_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_8_io_hostInterface_write_addr = io_hostInterface_8_write_addr; // @[CGRA.scala 595:36]
  assign lsus_8_io_hostInterface_write_data_valid = io_hostInterface_8_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_8_io_hostInterface_write_data_bits = io_hostInterface_8_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_8_io_hostInterface_cycle = io_hostInterface_8_cycle; // @[CGRA.scala 595:36]
  assign lsus_8_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_8_io_in_0 = gibs_16_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_8_io_in_1 = gibs_20_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_9_clock = clock;
  assign lsus_9_reset = reset;
  assign lsus_9_io_cfg_en = cfgRegs_10[46]; // @[CGRA.scala 678:35]
  assign lsus_9_io_cfg_addr = cfgRegs_10[45:32]; // @[CGRA.scala 679:37]
  assign lsus_9_io_cfg_data = cfgRegs_10[31:0]; // @[CGRA.scala 680:37]
  assign lsus_9_io_hostInterface_read_addr = io_hostInterface_9_read_addr; // @[CGRA.scala 595:36]
  assign lsus_9_io_hostInterface_read_data_ready = io_hostInterface_9_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_9_io_hostInterface_write_addr = io_hostInterface_9_write_addr; // @[CGRA.scala 595:36]
  assign lsus_9_io_hostInterface_write_data_valid = io_hostInterface_9_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_9_io_hostInterface_write_data_bits = io_hostInterface_9_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_9_io_hostInterface_cycle = io_hostInterface_9_cycle; // @[CGRA.scala 595:36]
  assign lsus_9_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_9_io_in_0 = gibs_19_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_9_io_in_1 = gibs_23_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_10_clock = clock;
  assign lsus_10_reset = reset;
  assign lsus_10_io_cfg_en = cfgRegs_12[46]; // @[CGRA.scala 678:35]
  assign lsus_10_io_cfg_addr = cfgRegs_12[45:32]; // @[CGRA.scala 679:37]
  assign lsus_10_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 680:37]
  assign lsus_10_io_hostInterface_read_addr = io_hostInterface_10_read_addr; // @[CGRA.scala 595:36]
  assign lsus_10_io_hostInterface_read_data_ready = io_hostInterface_10_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_10_io_hostInterface_write_addr = io_hostInterface_10_write_addr; // @[CGRA.scala 595:36]
  assign lsus_10_io_hostInterface_write_data_valid = io_hostInterface_10_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_10_io_hostInterface_write_data_bits = io_hostInterface_10_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_10_io_hostInterface_cycle = io_hostInterface_10_cycle; // @[CGRA.scala 595:36]
  assign lsus_10_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_10_io_in_0 = gibs_20_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_10_io_in_1 = gibs_24_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_11_clock = clock;
  assign lsus_11_reset = reset;
  assign lsus_11_io_cfg_en = cfgRegs_12[46]; // @[CGRA.scala 678:35]
  assign lsus_11_io_cfg_addr = cfgRegs_12[45:32]; // @[CGRA.scala 679:37]
  assign lsus_11_io_cfg_data = cfgRegs_12[31:0]; // @[CGRA.scala 680:37]
  assign lsus_11_io_hostInterface_read_addr = io_hostInterface_11_read_addr; // @[CGRA.scala 595:36]
  assign lsus_11_io_hostInterface_read_data_ready = io_hostInterface_11_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_11_io_hostInterface_write_addr = io_hostInterface_11_write_addr; // @[CGRA.scala 595:36]
  assign lsus_11_io_hostInterface_write_data_valid = io_hostInterface_11_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_11_io_hostInterface_write_data_bits = io_hostInterface_11_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_11_io_hostInterface_cycle = io_hostInterface_11_cycle; // @[CGRA.scala 595:36]
  assign lsus_11_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_11_io_in_0 = gibs_23_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_11_io_in_1 = gibs_27_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_12_clock = clock;
  assign lsus_12_reset = reset;
  assign lsus_12_io_cfg_en = cfgRegs_14[46]; // @[CGRA.scala 678:35]
  assign lsus_12_io_cfg_addr = cfgRegs_14[45:32]; // @[CGRA.scala 679:37]
  assign lsus_12_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 680:37]
  assign lsus_12_io_hostInterface_read_addr = io_hostInterface_12_read_addr; // @[CGRA.scala 595:36]
  assign lsus_12_io_hostInterface_read_data_ready = io_hostInterface_12_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_12_io_hostInterface_write_addr = io_hostInterface_12_write_addr; // @[CGRA.scala 595:36]
  assign lsus_12_io_hostInterface_write_data_valid = io_hostInterface_12_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_12_io_hostInterface_write_data_bits = io_hostInterface_12_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_12_io_hostInterface_cycle = io_hostInterface_12_cycle; // @[CGRA.scala 595:36]
  assign lsus_12_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_12_io_in_0 = gibs_24_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_12_io_in_1 = gibs_28_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_13_clock = clock;
  assign lsus_13_reset = reset;
  assign lsus_13_io_cfg_en = cfgRegs_14[46]; // @[CGRA.scala 678:35]
  assign lsus_13_io_cfg_addr = cfgRegs_14[45:32]; // @[CGRA.scala 679:37]
  assign lsus_13_io_cfg_data = cfgRegs_14[31:0]; // @[CGRA.scala 680:37]
  assign lsus_13_io_hostInterface_read_addr = io_hostInterface_13_read_addr; // @[CGRA.scala 595:36]
  assign lsus_13_io_hostInterface_read_data_ready = io_hostInterface_13_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_13_io_hostInterface_write_addr = io_hostInterface_13_write_addr; // @[CGRA.scala 595:36]
  assign lsus_13_io_hostInterface_write_data_valid = io_hostInterface_13_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_13_io_hostInterface_write_data_bits = io_hostInterface_13_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_13_io_hostInterface_cycle = io_hostInterface_13_cycle; // @[CGRA.scala 595:36]
  assign lsus_13_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_13_io_in_0 = gibs_27_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_13_io_in_1 = gibs_31_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_14_clock = clock;
  assign lsus_14_reset = reset;
  assign lsus_14_io_cfg_en = cfgRegs_16[46]; // @[CGRA.scala 678:35]
  assign lsus_14_io_cfg_addr = cfgRegs_16[45:32]; // @[CGRA.scala 679:37]
  assign lsus_14_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 680:37]
  assign lsus_14_io_hostInterface_read_addr = io_hostInterface_14_read_addr; // @[CGRA.scala 595:36]
  assign lsus_14_io_hostInterface_read_data_ready = io_hostInterface_14_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_14_io_hostInterface_write_addr = io_hostInterface_14_write_addr; // @[CGRA.scala 595:36]
  assign lsus_14_io_hostInterface_write_data_valid = io_hostInterface_14_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_14_io_hostInterface_write_data_bits = io_hostInterface_14_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_14_io_hostInterface_cycle = io_hostInterface_14_cycle; // @[CGRA.scala 595:36]
  assign lsus_14_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_14_io_in_0 = gibs_28_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_14_io_in_1 = gibs_32_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_15_clock = clock;
  assign lsus_15_reset = reset;
  assign lsus_15_io_cfg_en = cfgRegs_16[46]; // @[CGRA.scala 678:35]
  assign lsus_15_io_cfg_addr = cfgRegs_16[45:32]; // @[CGRA.scala 679:37]
  assign lsus_15_io_cfg_data = cfgRegs_16[31:0]; // @[CGRA.scala 680:37]
  assign lsus_15_io_hostInterface_read_addr = io_hostInterface_15_read_addr; // @[CGRA.scala 595:36]
  assign lsus_15_io_hostInterface_read_data_ready = io_hostInterface_15_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_15_io_hostInterface_write_addr = io_hostInterface_15_write_addr; // @[CGRA.scala 595:36]
  assign lsus_15_io_hostInterface_write_data_valid = io_hostInterface_15_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_15_io_hostInterface_write_data_bits = io_hostInterface_15_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_15_io_hostInterface_cycle = io_hostInterface_15_cycle; // @[CGRA.scala 595:36]
  assign lsus_15_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_15_io_in_0 = gibs_31_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_15_io_in_1 = gibs_35_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_16_clock = clock;
  assign lsus_16_reset = reset;
  assign lsus_16_io_cfg_en = cfgRegs_18[46]; // @[CGRA.scala 678:35]
  assign lsus_16_io_cfg_addr = cfgRegs_18[45:32]; // @[CGRA.scala 679:37]
  assign lsus_16_io_cfg_data = cfgRegs_18[31:0]; // @[CGRA.scala 680:37]
  assign lsus_16_io_hostInterface_read_addr = io_hostInterface_16_read_addr; // @[CGRA.scala 595:36]
  assign lsus_16_io_hostInterface_read_data_ready = io_hostInterface_16_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_16_io_hostInterface_write_addr = io_hostInterface_16_write_addr; // @[CGRA.scala 595:36]
  assign lsus_16_io_hostInterface_write_data_valid = io_hostInterface_16_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_16_io_hostInterface_write_data_bits = io_hostInterface_16_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_16_io_hostInterface_cycle = io_hostInterface_16_cycle; // @[CGRA.scala 595:36]
  assign lsus_16_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_16_io_in_0 = gibs_32_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_16_io_in_1 = gibs_36_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_17_clock = clock;
  assign lsus_17_reset = reset;
  assign lsus_17_io_cfg_en = cfgRegs_18[46]; // @[CGRA.scala 678:35]
  assign lsus_17_io_cfg_addr = cfgRegs_18[45:32]; // @[CGRA.scala 679:37]
  assign lsus_17_io_cfg_data = cfgRegs_18[31:0]; // @[CGRA.scala 680:37]
  assign lsus_17_io_hostInterface_read_addr = io_hostInterface_17_read_addr; // @[CGRA.scala 595:36]
  assign lsus_17_io_hostInterface_read_data_ready = io_hostInterface_17_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_17_io_hostInterface_write_addr = io_hostInterface_17_write_addr; // @[CGRA.scala 595:36]
  assign lsus_17_io_hostInterface_write_data_valid = io_hostInterface_17_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_17_io_hostInterface_write_data_bits = io_hostInterface_17_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_17_io_hostInterface_cycle = io_hostInterface_17_cycle; // @[CGRA.scala 595:36]
  assign lsus_17_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_17_io_in_0 = gibs_35_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_17_io_in_1 = gibs_39_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_18_clock = clock;
  assign lsus_18_reset = reset;
  assign lsus_18_io_cfg_en = cfgRegs_20[46]; // @[CGRA.scala 678:35]
  assign lsus_18_io_cfg_addr = cfgRegs_20[45:32]; // @[CGRA.scala 679:37]
  assign lsus_18_io_cfg_data = cfgRegs_20[31:0]; // @[CGRA.scala 680:37]
  assign lsus_18_io_hostInterface_read_addr = io_hostInterface_18_read_addr; // @[CGRA.scala 595:36]
  assign lsus_18_io_hostInterface_read_data_ready = io_hostInterface_18_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_18_io_hostInterface_write_addr = io_hostInterface_18_write_addr; // @[CGRA.scala 595:36]
  assign lsus_18_io_hostInterface_write_data_valid = io_hostInterface_18_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_18_io_hostInterface_write_data_bits = io_hostInterface_18_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_18_io_hostInterface_cycle = io_hostInterface_18_cycle; // @[CGRA.scala 595:36]
  assign lsus_18_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_18_io_in_0 = gibs_36_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_18_io_in_1 = gibs_40_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_19_clock = clock;
  assign lsus_19_reset = reset;
  assign lsus_19_io_cfg_en = cfgRegs_20[46]; // @[CGRA.scala 678:35]
  assign lsus_19_io_cfg_addr = cfgRegs_20[45:32]; // @[CGRA.scala 679:37]
  assign lsus_19_io_cfg_data = cfgRegs_20[31:0]; // @[CGRA.scala 680:37]
  assign lsus_19_io_hostInterface_read_addr = io_hostInterface_19_read_addr; // @[CGRA.scala 595:36]
  assign lsus_19_io_hostInterface_read_data_ready = io_hostInterface_19_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_19_io_hostInterface_write_addr = io_hostInterface_19_write_addr; // @[CGRA.scala 595:36]
  assign lsus_19_io_hostInterface_write_data_valid = io_hostInterface_19_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_19_io_hostInterface_write_data_bits = io_hostInterface_19_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_19_io_hostInterface_cycle = io_hostInterface_19_cycle; // @[CGRA.scala 595:36]
  assign lsus_19_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_19_io_in_0 = gibs_39_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_19_io_in_1 = gibs_43_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_20_clock = clock;
  assign lsus_20_reset = reset;
  assign lsus_20_io_cfg_en = cfgRegs_22[46]; // @[CGRA.scala 678:35]
  assign lsus_20_io_cfg_addr = cfgRegs_22[45:32]; // @[CGRA.scala 679:37]
  assign lsus_20_io_cfg_data = cfgRegs_22[31:0]; // @[CGRA.scala 680:37]
  assign lsus_20_io_hostInterface_read_addr = io_hostInterface_20_read_addr; // @[CGRA.scala 595:36]
  assign lsus_20_io_hostInterface_read_data_ready = io_hostInterface_20_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_20_io_hostInterface_write_addr = io_hostInterface_20_write_addr; // @[CGRA.scala 595:36]
  assign lsus_20_io_hostInterface_write_data_valid = io_hostInterface_20_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_20_io_hostInterface_write_data_bits = io_hostInterface_20_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_20_io_hostInterface_cycle = io_hostInterface_20_cycle; // @[CGRA.scala 595:36]
  assign lsus_20_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_20_io_in_0 = gibs_40_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_20_io_in_1 = gibs_44_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_21_clock = clock;
  assign lsus_21_reset = reset;
  assign lsus_21_io_cfg_en = cfgRegs_22[46]; // @[CGRA.scala 678:35]
  assign lsus_21_io_cfg_addr = cfgRegs_22[45:32]; // @[CGRA.scala 679:37]
  assign lsus_21_io_cfg_data = cfgRegs_22[31:0]; // @[CGRA.scala 680:37]
  assign lsus_21_io_hostInterface_read_addr = io_hostInterface_21_read_addr; // @[CGRA.scala 595:36]
  assign lsus_21_io_hostInterface_read_data_ready = io_hostInterface_21_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_21_io_hostInterface_write_addr = io_hostInterface_21_write_addr; // @[CGRA.scala 595:36]
  assign lsus_21_io_hostInterface_write_data_valid = io_hostInterface_21_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_21_io_hostInterface_write_data_bits = io_hostInterface_21_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_21_io_hostInterface_cycle = io_hostInterface_21_cycle; // @[CGRA.scala 595:36]
  assign lsus_21_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_21_io_in_0 = gibs_43_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_21_io_in_1 = gibs_47_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_22_clock = clock;
  assign lsus_22_reset = reset;
  assign lsus_22_io_cfg_en = cfgRegs_24[46]; // @[CGRA.scala 678:35]
  assign lsus_22_io_cfg_addr = cfgRegs_24[45:32]; // @[CGRA.scala 679:37]
  assign lsus_22_io_cfg_data = cfgRegs_24[31:0]; // @[CGRA.scala 680:37]
  assign lsus_22_io_hostInterface_read_addr = io_hostInterface_22_read_addr; // @[CGRA.scala 595:36]
  assign lsus_22_io_hostInterface_read_data_ready = io_hostInterface_22_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_22_io_hostInterface_write_addr = io_hostInterface_22_write_addr; // @[CGRA.scala 595:36]
  assign lsus_22_io_hostInterface_write_data_valid = io_hostInterface_22_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_22_io_hostInterface_write_data_bits = io_hostInterface_22_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_22_io_hostInterface_cycle = io_hostInterface_22_cycle; // @[CGRA.scala 595:36]
  assign lsus_22_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_22_io_in_0 = gibs_44_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_22_io_in_1 = gibs_48_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_23_clock = clock;
  assign lsus_23_reset = reset;
  assign lsus_23_io_cfg_en = cfgRegs_24[46]; // @[CGRA.scala 678:35]
  assign lsus_23_io_cfg_addr = cfgRegs_24[45:32]; // @[CGRA.scala 679:37]
  assign lsus_23_io_cfg_data = cfgRegs_24[31:0]; // @[CGRA.scala 680:37]
  assign lsus_23_io_hostInterface_read_addr = io_hostInterface_23_read_addr; // @[CGRA.scala 595:36]
  assign lsus_23_io_hostInterface_read_data_ready = io_hostInterface_23_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_23_io_hostInterface_write_addr = io_hostInterface_23_write_addr; // @[CGRA.scala 595:36]
  assign lsus_23_io_hostInterface_write_data_valid = io_hostInterface_23_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_23_io_hostInterface_write_data_bits = io_hostInterface_23_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_23_io_hostInterface_cycle = io_hostInterface_23_cycle; // @[CGRA.scala 595:36]
  assign lsus_23_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_23_io_in_0 = gibs_47_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_23_io_in_1 = gibs_51_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_24_clock = clock;
  assign lsus_24_reset = reset;
  assign lsus_24_io_cfg_en = cfgRegs_26[46]; // @[CGRA.scala 678:35]
  assign lsus_24_io_cfg_addr = cfgRegs_26[45:32]; // @[CGRA.scala 679:37]
  assign lsus_24_io_cfg_data = cfgRegs_26[31:0]; // @[CGRA.scala 680:37]
  assign lsus_24_io_hostInterface_read_addr = io_hostInterface_24_read_addr; // @[CGRA.scala 595:36]
  assign lsus_24_io_hostInterface_read_data_ready = io_hostInterface_24_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_24_io_hostInterface_write_addr = io_hostInterface_24_write_addr; // @[CGRA.scala 595:36]
  assign lsus_24_io_hostInterface_write_data_valid = io_hostInterface_24_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_24_io_hostInterface_write_data_bits = io_hostInterface_24_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_24_io_hostInterface_cycle = io_hostInterface_24_cycle; // @[CGRA.scala 595:36]
  assign lsus_24_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_24_io_in_0 = gibs_48_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_24_io_in_1 = gibs_52_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_25_clock = clock;
  assign lsus_25_reset = reset;
  assign lsus_25_io_cfg_en = cfgRegs_26[46]; // @[CGRA.scala 678:35]
  assign lsus_25_io_cfg_addr = cfgRegs_26[45:32]; // @[CGRA.scala 679:37]
  assign lsus_25_io_cfg_data = cfgRegs_26[31:0]; // @[CGRA.scala 680:37]
  assign lsus_25_io_hostInterface_read_addr = io_hostInterface_25_read_addr; // @[CGRA.scala 595:36]
  assign lsus_25_io_hostInterface_read_data_ready = io_hostInterface_25_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_25_io_hostInterface_write_addr = io_hostInterface_25_write_addr; // @[CGRA.scala 595:36]
  assign lsus_25_io_hostInterface_write_data_valid = io_hostInterface_25_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_25_io_hostInterface_write_data_bits = io_hostInterface_25_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_25_io_hostInterface_cycle = io_hostInterface_25_cycle; // @[CGRA.scala 595:36]
  assign lsus_25_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_25_io_in_0 = gibs_51_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_25_io_in_1 = gibs_55_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_26_clock = clock;
  assign lsus_26_reset = reset;
  assign lsus_26_io_cfg_en = cfgRegs_28[46]; // @[CGRA.scala 678:35]
  assign lsus_26_io_cfg_addr = cfgRegs_28[45:32]; // @[CGRA.scala 679:37]
  assign lsus_26_io_cfg_data = cfgRegs_28[31:0]; // @[CGRA.scala 680:37]
  assign lsus_26_io_hostInterface_read_addr = io_hostInterface_26_read_addr; // @[CGRA.scala 595:36]
  assign lsus_26_io_hostInterface_read_data_ready = io_hostInterface_26_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_26_io_hostInterface_write_addr = io_hostInterface_26_write_addr; // @[CGRA.scala 595:36]
  assign lsus_26_io_hostInterface_write_data_valid = io_hostInterface_26_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_26_io_hostInterface_write_data_bits = io_hostInterface_26_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_26_io_hostInterface_cycle = io_hostInterface_26_cycle; // @[CGRA.scala 595:36]
  assign lsus_26_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_26_io_in_0 = gibs_52_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_26_io_in_1 = gibs_56_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_27_clock = clock;
  assign lsus_27_reset = reset;
  assign lsus_27_io_cfg_en = cfgRegs_28[46]; // @[CGRA.scala 678:35]
  assign lsus_27_io_cfg_addr = cfgRegs_28[45:32]; // @[CGRA.scala 679:37]
  assign lsus_27_io_cfg_data = cfgRegs_28[31:0]; // @[CGRA.scala 680:37]
  assign lsus_27_io_hostInterface_read_addr = io_hostInterface_27_read_addr; // @[CGRA.scala 595:36]
  assign lsus_27_io_hostInterface_read_data_ready = io_hostInterface_27_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_27_io_hostInterface_write_addr = io_hostInterface_27_write_addr; // @[CGRA.scala 595:36]
  assign lsus_27_io_hostInterface_write_data_valid = io_hostInterface_27_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_27_io_hostInterface_write_data_bits = io_hostInterface_27_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_27_io_hostInterface_cycle = io_hostInterface_27_cycle; // @[CGRA.scala 595:36]
  assign lsus_27_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_27_io_in_0 = gibs_55_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_27_io_in_1 = gibs_59_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_28_clock = clock;
  assign lsus_28_reset = reset;
  assign lsus_28_io_cfg_en = cfgRegs_30[46]; // @[CGRA.scala 678:35]
  assign lsus_28_io_cfg_addr = cfgRegs_30[45:32]; // @[CGRA.scala 679:37]
  assign lsus_28_io_cfg_data = cfgRegs_30[31:0]; // @[CGRA.scala 680:37]
  assign lsus_28_io_hostInterface_read_addr = io_hostInterface_28_read_addr; // @[CGRA.scala 595:36]
  assign lsus_28_io_hostInterface_read_data_ready = io_hostInterface_28_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_28_io_hostInterface_write_addr = io_hostInterface_28_write_addr; // @[CGRA.scala 595:36]
  assign lsus_28_io_hostInterface_write_data_valid = io_hostInterface_28_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_28_io_hostInterface_write_data_bits = io_hostInterface_28_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_28_io_hostInterface_cycle = io_hostInterface_28_cycle; // @[CGRA.scala 595:36]
  assign lsus_28_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_28_io_in_0 = gibs_56_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_28_io_in_1 = gibs_60_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_29_clock = clock;
  assign lsus_29_reset = reset;
  assign lsus_29_io_cfg_en = cfgRegs_30[46]; // @[CGRA.scala 678:35]
  assign lsus_29_io_cfg_addr = cfgRegs_30[45:32]; // @[CGRA.scala 679:37]
  assign lsus_29_io_cfg_data = cfgRegs_30[31:0]; // @[CGRA.scala 680:37]
  assign lsus_29_io_hostInterface_read_addr = io_hostInterface_29_read_addr; // @[CGRA.scala 595:36]
  assign lsus_29_io_hostInterface_read_data_ready = io_hostInterface_29_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_29_io_hostInterface_write_addr = io_hostInterface_29_write_addr; // @[CGRA.scala 595:36]
  assign lsus_29_io_hostInterface_write_data_valid = io_hostInterface_29_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_29_io_hostInterface_write_data_bits = io_hostInterface_29_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_29_io_hostInterface_cycle = io_hostInterface_29_cycle; // @[CGRA.scala 595:36]
  assign lsus_29_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_29_io_in_0 = gibs_59_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_29_io_in_1 = gibs_63_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_30_clock = clock;
  assign lsus_30_reset = reset;
  assign lsus_30_io_cfg_en = cfgRegs_32[46]; // @[CGRA.scala 678:35]
  assign lsus_30_io_cfg_addr = cfgRegs_32[45:32]; // @[CGRA.scala 679:37]
  assign lsus_30_io_cfg_data = cfgRegs_32[31:0]; // @[CGRA.scala 680:37]
  assign lsus_30_io_hostInterface_read_addr = io_hostInterface_30_read_addr; // @[CGRA.scala 595:36]
  assign lsus_30_io_hostInterface_read_data_ready = io_hostInterface_30_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_30_io_hostInterface_write_addr = io_hostInterface_30_write_addr; // @[CGRA.scala 595:36]
  assign lsus_30_io_hostInterface_write_data_valid = io_hostInterface_30_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_30_io_hostInterface_write_data_bits = io_hostInterface_30_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_30_io_hostInterface_cycle = io_hostInterface_30_cycle; // @[CGRA.scala 595:36]
  assign lsus_30_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_30_io_in_0 = gibs_60_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_30_io_in_1 = gibs_64_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_31_clock = clock;
  assign lsus_31_reset = reset;
  assign lsus_31_io_cfg_en = cfgRegs_32[46]; // @[CGRA.scala 678:35]
  assign lsus_31_io_cfg_addr = cfgRegs_32[45:32]; // @[CGRA.scala 679:37]
  assign lsus_31_io_cfg_data = cfgRegs_32[31:0]; // @[CGRA.scala 680:37]
  assign lsus_31_io_hostInterface_read_addr = io_hostInterface_31_read_addr; // @[CGRA.scala 595:36]
  assign lsus_31_io_hostInterface_read_data_ready = io_hostInterface_31_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_31_io_hostInterface_write_addr = io_hostInterface_31_write_addr; // @[CGRA.scala 595:36]
  assign lsus_31_io_hostInterface_write_data_valid = io_hostInterface_31_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_31_io_hostInterface_write_data_bits = io_hostInterface_31_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_31_io_hostInterface_cycle = io_hostInterface_31_cycle; // @[CGRA.scala 595:36]
  assign lsus_31_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_31_io_in_0 = gibs_63_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_31_io_in_1 = gibs_67_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_32_clock = clock;
  assign lsus_32_reset = reset;
  assign lsus_32_io_cfg_en = cfgRegs_34[46]; // @[CGRA.scala 678:35]
  assign lsus_32_io_cfg_addr = cfgRegs_34[45:32]; // @[CGRA.scala 679:37]
  assign lsus_32_io_cfg_data = cfgRegs_34[31:0]; // @[CGRA.scala 680:37]
  assign lsus_32_io_hostInterface_read_addr = io_hostInterface_32_read_addr; // @[CGRA.scala 595:36]
  assign lsus_32_io_hostInterface_read_data_ready = io_hostInterface_32_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_32_io_hostInterface_write_addr = io_hostInterface_32_write_addr; // @[CGRA.scala 595:36]
  assign lsus_32_io_hostInterface_write_data_valid = io_hostInterface_32_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_32_io_hostInterface_write_data_bits = io_hostInterface_32_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_32_io_hostInterface_cycle = io_hostInterface_32_cycle; // @[CGRA.scala 595:36]
  assign lsus_32_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_32_io_in_0 = gibs_64_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_32_io_in_1 = gibs_68_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_33_clock = clock;
  assign lsus_33_reset = reset;
  assign lsus_33_io_cfg_en = cfgRegs_34[46]; // @[CGRA.scala 678:35]
  assign lsus_33_io_cfg_addr = cfgRegs_34[45:32]; // @[CGRA.scala 679:37]
  assign lsus_33_io_cfg_data = cfgRegs_34[31:0]; // @[CGRA.scala 680:37]
  assign lsus_33_io_hostInterface_read_addr = io_hostInterface_33_read_addr; // @[CGRA.scala 595:36]
  assign lsus_33_io_hostInterface_read_data_ready = io_hostInterface_33_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_33_io_hostInterface_write_addr = io_hostInterface_33_write_addr; // @[CGRA.scala 595:36]
  assign lsus_33_io_hostInterface_write_data_valid = io_hostInterface_33_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_33_io_hostInterface_write_data_bits = io_hostInterface_33_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_33_io_hostInterface_cycle = io_hostInterface_33_cycle; // @[CGRA.scala 595:36]
  assign lsus_33_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_33_io_in_0 = gibs_67_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_33_io_in_1 = gibs_71_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_34_clock = clock;
  assign lsus_34_reset = reset;
  assign lsus_34_io_cfg_en = cfgRegs_36[46]; // @[CGRA.scala 678:35]
  assign lsus_34_io_cfg_addr = cfgRegs_36[45:32]; // @[CGRA.scala 679:37]
  assign lsus_34_io_cfg_data = cfgRegs_36[31:0]; // @[CGRA.scala 680:37]
  assign lsus_34_io_hostInterface_read_addr = io_hostInterface_34_read_addr; // @[CGRA.scala 595:36]
  assign lsus_34_io_hostInterface_read_data_ready = io_hostInterface_34_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_34_io_hostInterface_write_addr = io_hostInterface_34_write_addr; // @[CGRA.scala 595:36]
  assign lsus_34_io_hostInterface_write_data_valid = io_hostInterface_34_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_34_io_hostInterface_write_data_bits = io_hostInterface_34_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_34_io_hostInterface_cycle = io_hostInterface_34_cycle; // @[CGRA.scala 595:36]
  assign lsus_34_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_34_io_in_0 = gibs_68_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_34_io_in_1 = gibs_72_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_35_clock = clock;
  assign lsus_35_reset = reset;
  assign lsus_35_io_cfg_en = cfgRegs_36[46]; // @[CGRA.scala 678:35]
  assign lsus_35_io_cfg_addr = cfgRegs_36[45:32]; // @[CGRA.scala 679:37]
  assign lsus_35_io_cfg_data = cfgRegs_36[31:0]; // @[CGRA.scala 680:37]
  assign lsus_35_io_hostInterface_read_addr = io_hostInterface_35_read_addr; // @[CGRA.scala 595:36]
  assign lsus_35_io_hostInterface_read_data_ready = io_hostInterface_35_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_35_io_hostInterface_write_addr = io_hostInterface_35_write_addr; // @[CGRA.scala 595:36]
  assign lsus_35_io_hostInterface_write_data_valid = io_hostInterface_35_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_35_io_hostInterface_write_data_bits = io_hostInterface_35_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_35_io_hostInterface_cycle = io_hostInterface_35_cycle; // @[CGRA.scala 595:36]
  assign lsus_35_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_35_io_in_0 = gibs_71_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_35_io_in_1 = gibs_75_io_ipinNE_0; // @[CGRA.scala 623:16]
  assign lsus_36_clock = clock;
  assign lsus_36_reset = reset;
  assign lsus_36_io_cfg_en = cfgRegs_38[46]; // @[CGRA.scala 678:35]
  assign lsus_36_io_cfg_addr = cfgRegs_38[45:32]; // @[CGRA.scala 679:37]
  assign lsus_36_io_cfg_data = cfgRegs_38[31:0]; // @[CGRA.scala 680:37]
  assign lsus_36_io_hostInterface_read_addr = io_hostInterface_36_read_addr; // @[CGRA.scala 595:36]
  assign lsus_36_io_hostInterface_read_data_ready = io_hostInterface_36_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_36_io_hostInterface_write_addr = io_hostInterface_36_write_addr; // @[CGRA.scala 595:36]
  assign lsus_36_io_hostInterface_write_data_valid = io_hostInterface_36_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_36_io_hostInterface_write_data_bits = io_hostInterface_36_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_36_io_hostInterface_cycle = io_hostInterface_36_cycle; // @[CGRA.scala 595:36]
  assign lsus_36_io_en = io_en_0; // @[CGRA.scala 594:25]
  assign lsus_36_io_in_0 = gibs_72_io_ipinSW_0; // @[CGRA.scala 599:14]
  assign lsus_36_io_in_1 = gibs_76_io_ipinNW_0; // @[CGRA.scala 603:14]
  assign lsus_37_clock = clock;
  assign lsus_37_reset = reset;
  assign lsus_37_io_cfg_en = cfgRegs_38[46]; // @[CGRA.scala 678:35]
  assign lsus_37_io_cfg_addr = cfgRegs_38[45:32]; // @[CGRA.scala 679:37]
  assign lsus_37_io_cfg_data = cfgRegs_38[31:0]; // @[CGRA.scala 680:37]
  assign lsus_37_io_hostInterface_read_addr = io_hostInterface_37_read_addr; // @[CGRA.scala 595:36]
  assign lsus_37_io_hostInterface_read_data_ready = io_hostInterface_37_read_data_ready; // @[CGRA.scala 595:36]
  assign lsus_37_io_hostInterface_write_addr = io_hostInterface_37_write_addr; // @[CGRA.scala 595:36]
  assign lsus_37_io_hostInterface_write_data_valid = io_hostInterface_37_write_data_valid; // @[CGRA.scala 595:36]
  assign lsus_37_io_hostInterface_write_data_bits = io_hostInterface_37_write_data_bits; // @[CGRA.scala 595:36]
  assign lsus_37_io_hostInterface_cycle = io_hostInterface_37_cycle; // @[CGRA.scala 595:36]
  assign lsus_37_io_en = io_en_4; // @[CGRA.scala 594:25]
  assign lsus_37_io_in_0 = gibs_75_io_ipinSE_0; // @[CGRA.scala 619:16]
  assign lsus_37_io_in_1 = gibs_79_io_ipinNE_0; // @[CGRA.scala 623:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cfgRegs_0 = _RAND_0[46:0];
  _RAND_1 = {2{`RANDOM}};
  cfgRegs_1 = _RAND_1[46:0];
  _RAND_2 = {2{`RANDOM}};
  cfgRegs_2 = _RAND_2[46:0];
  _RAND_3 = {2{`RANDOM}};
  cfgRegs_3 = _RAND_3[46:0];
  _RAND_4 = {2{`RANDOM}};
  cfgRegs_4 = _RAND_4[46:0];
  _RAND_5 = {2{`RANDOM}};
  cfgRegs_5 = _RAND_5[46:0];
  _RAND_6 = {2{`RANDOM}};
  cfgRegs_6 = _RAND_6[46:0];
  _RAND_7 = {2{`RANDOM}};
  cfgRegs_7 = _RAND_7[46:0];
  _RAND_8 = {2{`RANDOM}};
  cfgRegs_8 = _RAND_8[46:0];
  _RAND_9 = {2{`RANDOM}};
  cfgRegs_9 = _RAND_9[46:0];
  _RAND_10 = {2{`RANDOM}};
  cfgRegs_10 = _RAND_10[46:0];
  _RAND_11 = {2{`RANDOM}};
  cfgRegs_11 = _RAND_11[46:0];
  _RAND_12 = {2{`RANDOM}};
  cfgRegs_12 = _RAND_12[46:0];
  _RAND_13 = {2{`RANDOM}};
  cfgRegs_13 = _RAND_13[46:0];
  _RAND_14 = {2{`RANDOM}};
  cfgRegs_14 = _RAND_14[46:0];
  _RAND_15 = {2{`RANDOM}};
  cfgRegs_15 = _RAND_15[46:0];
  _RAND_16 = {2{`RANDOM}};
  cfgRegs_16 = _RAND_16[46:0];
  _RAND_17 = {2{`RANDOM}};
  cfgRegs_17 = _RAND_17[46:0];
  _RAND_18 = {2{`RANDOM}};
  cfgRegs_18 = _RAND_18[46:0];
  _RAND_19 = {2{`RANDOM}};
  cfgRegs_19 = _RAND_19[46:0];
  _RAND_20 = {2{`RANDOM}};
  cfgRegs_20 = _RAND_20[46:0];
  _RAND_21 = {2{`RANDOM}};
  cfgRegs_21 = _RAND_21[46:0];
  _RAND_22 = {2{`RANDOM}};
  cfgRegs_22 = _RAND_22[46:0];
  _RAND_23 = {2{`RANDOM}};
  cfgRegs_23 = _RAND_23[46:0];
  _RAND_24 = {2{`RANDOM}};
  cfgRegs_24 = _RAND_24[46:0];
  _RAND_25 = {2{`RANDOM}};
  cfgRegs_25 = _RAND_25[46:0];
  _RAND_26 = {2{`RANDOM}};
  cfgRegs_26 = _RAND_26[46:0];
  _RAND_27 = {2{`RANDOM}};
  cfgRegs_27 = _RAND_27[46:0];
  _RAND_28 = {2{`RANDOM}};
  cfgRegs_28 = _RAND_28[46:0];
  _RAND_29 = {2{`RANDOM}};
  cfgRegs_29 = _RAND_29[46:0];
  _RAND_30 = {2{`RANDOM}};
  cfgRegs_30 = _RAND_30[46:0];
  _RAND_31 = {2{`RANDOM}};
  cfgRegs_31 = _RAND_31[46:0];
  _RAND_32 = {2{`RANDOM}};
  cfgRegs_32 = _RAND_32[46:0];
  _RAND_33 = {2{`RANDOM}};
  cfgRegs_33 = _RAND_33[46:0];
  _RAND_34 = {2{`RANDOM}};
  cfgRegs_34 = _RAND_34[46:0];
  _RAND_35 = {2{`RANDOM}};
  cfgRegs_35 = _RAND_35[46:0];
  _RAND_36 = {2{`RANDOM}};
  cfgRegs_36 = _RAND_36[46:0];
  _RAND_37 = {2{`RANDOM}};
  cfgRegs_37 = _RAND_37[46:0];
  _RAND_38 = {2{`RANDOM}};
  cfgRegs_38 = _RAND_38[46:0];
  _RAND_39 = {2{`RANDOM}};
  cfgRegs_39 = _RAND_39[46:0];
  _RAND_40 = {2{`RANDOM}};
  cfgRegs_40 = _RAND_40[46:0];
  _RAND_41 = {2{`RANDOM}};
  cfgRegs_41 = _RAND_41[46:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cfgRegs_0 <= 47'h0;
    end else begin
      cfgRegs_0 <= _T_2;
    end
    if (reset) begin
      cfgRegs_1 <= 47'h0;
    end else begin
      cfgRegs_1 <= cfgRegs_0;
    end
    if (reset) begin
      cfgRegs_2 <= 47'h0;
    end else begin
      cfgRegs_2 <= cfgRegs_1;
    end
    if (reset) begin
      cfgRegs_3 <= 47'h0;
    end else begin
      cfgRegs_3 <= cfgRegs_2;
    end
    if (reset) begin
      cfgRegs_4 <= 47'h0;
    end else begin
      cfgRegs_4 <= cfgRegs_3;
    end
    if (reset) begin
      cfgRegs_5 <= 47'h0;
    end else begin
      cfgRegs_5 <= cfgRegs_4;
    end
    if (reset) begin
      cfgRegs_6 <= 47'h0;
    end else begin
      cfgRegs_6 <= cfgRegs_5;
    end
    if (reset) begin
      cfgRegs_7 <= 47'h0;
    end else begin
      cfgRegs_7 <= cfgRegs_6;
    end
    if (reset) begin
      cfgRegs_8 <= 47'h0;
    end else begin
      cfgRegs_8 <= cfgRegs_7;
    end
    if (reset) begin
      cfgRegs_9 <= 47'h0;
    end else begin
      cfgRegs_9 <= cfgRegs_8;
    end
    if (reset) begin
      cfgRegs_10 <= 47'h0;
    end else begin
      cfgRegs_10 <= cfgRegs_9;
    end
    if (reset) begin
      cfgRegs_11 <= 47'h0;
    end else begin
      cfgRegs_11 <= cfgRegs_10;
    end
    if (reset) begin
      cfgRegs_12 <= 47'h0;
    end else begin
      cfgRegs_12 <= cfgRegs_11;
    end
    if (reset) begin
      cfgRegs_13 <= 47'h0;
    end else begin
      cfgRegs_13 <= cfgRegs_12;
    end
    if (reset) begin
      cfgRegs_14 <= 47'h0;
    end else begin
      cfgRegs_14 <= cfgRegs_13;
    end
    if (reset) begin
      cfgRegs_15 <= 47'h0;
    end else begin
      cfgRegs_15 <= cfgRegs_14;
    end
    if (reset) begin
      cfgRegs_16 <= 47'h0;
    end else begin
      cfgRegs_16 <= cfgRegs_15;
    end
    if (reset) begin
      cfgRegs_17 <= 47'h0;
    end else begin
      cfgRegs_17 <= cfgRegs_16;
    end
    if (reset) begin
      cfgRegs_18 <= 47'h0;
    end else begin
      cfgRegs_18 <= cfgRegs_17;
    end
    if (reset) begin
      cfgRegs_19 <= 47'h0;
    end else begin
      cfgRegs_19 <= cfgRegs_18;
    end
    if (reset) begin
      cfgRegs_20 <= 47'h0;
    end else begin
      cfgRegs_20 <= cfgRegs_19;
    end
    if (reset) begin
      cfgRegs_21 <= 47'h0;
    end else begin
      cfgRegs_21 <= cfgRegs_20;
    end
    if (reset) begin
      cfgRegs_22 <= 47'h0;
    end else begin
      cfgRegs_22 <= cfgRegs_21;
    end
    if (reset) begin
      cfgRegs_23 <= 47'h0;
    end else begin
      cfgRegs_23 <= cfgRegs_22;
    end
    if (reset) begin
      cfgRegs_24 <= 47'h0;
    end else begin
      cfgRegs_24 <= cfgRegs_23;
    end
    if (reset) begin
      cfgRegs_25 <= 47'h0;
    end else begin
      cfgRegs_25 <= cfgRegs_24;
    end
    if (reset) begin
      cfgRegs_26 <= 47'h0;
    end else begin
      cfgRegs_26 <= cfgRegs_25;
    end
    if (reset) begin
      cfgRegs_27 <= 47'h0;
    end else begin
      cfgRegs_27 <= cfgRegs_26;
    end
    if (reset) begin
      cfgRegs_28 <= 47'h0;
    end else begin
      cfgRegs_28 <= cfgRegs_27;
    end
    if (reset) begin
      cfgRegs_29 <= 47'h0;
    end else begin
      cfgRegs_29 <= cfgRegs_28;
    end
    if (reset) begin
      cfgRegs_30 <= 47'h0;
    end else begin
      cfgRegs_30 <= cfgRegs_29;
    end
    if (reset) begin
      cfgRegs_31 <= 47'h0;
    end else begin
      cfgRegs_31 <= cfgRegs_30;
    end
    if (reset) begin
      cfgRegs_32 <= 47'h0;
    end else begin
      cfgRegs_32 <= cfgRegs_31;
    end
    if (reset) begin
      cfgRegs_33 <= 47'h0;
    end else begin
      cfgRegs_33 <= cfgRegs_32;
    end
    if (reset) begin
      cfgRegs_34 <= 47'h0;
    end else begin
      cfgRegs_34 <= cfgRegs_33;
    end
    if (reset) begin
      cfgRegs_35 <= 47'h0;
    end else begin
      cfgRegs_35 <= cfgRegs_34;
    end
    if (reset) begin
      cfgRegs_36 <= 47'h0;
    end else begin
      cfgRegs_36 <= cfgRegs_35;
    end
    if (reset) begin
      cfgRegs_37 <= 47'h0;
    end else begin
      cfgRegs_37 <= cfgRegs_36;
    end
    if (reset) begin
      cfgRegs_38 <= 47'h0;
    end else begin
      cfgRegs_38 <= cfgRegs_37;
    end
    if (reset) begin
      cfgRegs_39 <= 47'h0;
    end else begin
      cfgRegs_39 <= cfgRegs_38;
    end
    if (reset) begin
      cfgRegs_40 <= 47'h0;
    end else begin
      cfgRegs_40 <= cfgRegs_39;
    end
    if (reset) begin
      cfgRegs_41 <= 47'h0;
    end else begin
      cfgRegs_41 <= cfgRegs_40;
    end
  end
endmodule
