module Dispatch(
  input  [1151:0] io_configuration,
  output [5:0]    io_outs_191,
  output [5:0]    io_outs_190,
  output [5:0]    io_outs_189,
  output [5:0]    io_outs_188,
  output [5:0]    io_outs_187,
  output [5:0]    io_outs_186,
  output [5:0]    io_outs_185,
  output [5:0]    io_outs_184,
  output [5:0]    io_outs_183,
  output [5:0]    io_outs_182,
  output [5:0]    io_outs_181,
  output [5:0]    io_outs_180,
  output [5:0]    io_outs_179,
  output [5:0]    io_outs_178,
  output [5:0]    io_outs_177,
  output [5:0]    io_outs_176,
  output [5:0]    io_outs_175,
  output [5:0]    io_outs_174,
  output [5:0]    io_outs_173,
  output [5:0]    io_outs_172,
  output [5:0]    io_outs_171,
  output [5:0]    io_outs_170,
  output [5:0]    io_outs_169,
  output [5:0]    io_outs_168,
  output [5:0]    io_outs_167,
  output [5:0]    io_outs_166,
  output [5:0]    io_outs_165,
  output [5:0]    io_outs_164,
  output [5:0]    io_outs_163,
  output [5:0]    io_outs_162,
  output [5:0]    io_outs_161,
  output [5:0]    io_outs_160,
  output [5:0]    io_outs_159,
  output [5:0]    io_outs_158,
  output [5:0]    io_outs_157,
  output [5:0]    io_outs_156,
  output [5:0]    io_outs_155,
  output [5:0]    io_outs_154,
  output [5:0]    io_outs_153,
  output [5:0]    io_outs_152,
  output [5:0]    io_outs_151,
  output [5:0]    io_outs_150,
  output [5:0]    io_outs_149,
  output [5:0]    io_outs_148,
  output [5:0]    io_outs_147,
  output [5:0]    io_outs_146,
  output [5:0]    io_outs_145,
  output [5:0]    io_outs_144,
  output [5:0]    io_outs_143,
  output [5:0]    io_outs_142,
  output [5:0]    io_outs_141,
  output [5:0]    io_outs_140,
  output [5:0]    io_outs_139,
  output [5:0]    io_outs_138,
  output [5:0]    io_outs_137,
  output [5:0]    io_outs_136,
  output [5:0]    io_outs_135,
  output [5:0]    io_outs_134,
  output [5:0]    io_outs_133,
  output [5:0]    io_outs_132,
  output [5:0]    io_outs_131,
  output [5:0]    io_outs_130,
  output [5:0]    io_outs_129,
  output [5:0]    io_outs_128,
  output [5:0]    io_outs_127,
  output [5:0]    io_outs_126,
  output [5:0]    io_outs_125,
  output [5:0]    io_outs_124,
  output [5:0]    io_outs_123,
  output [5:0]    io_outs_122,
  output [5:0]    io_outs_121,
  output [5:0]    io_outs_120,
  output [5:0]    io_outs_119,
  output [5:0]    io_outs_118,
  output [5:0]    io_outs_117,
  output [5:0]    io_outs_116,
  output [5:0]    io_outs_115,
  output [5:0]    io_outs_114,
  output [5:0]    io_outs_113,
  output [5:0]    io_outs_112,
  output [5:0]    io_outs_111,
  output [5:0]    io_outs_110,
  output [5:0]    io_outs_109,
  output [5:0]    io_outs_108,
  output [5:0]    io_outs_107,
  output [5:0]    io_outs_106,
  output [5:0]    io_outs_105,
  output [5:0]    io_outs_104,
  output [5:0]    io_outs_103,
  output [5:0]    io_outs_102,
  output [5:0]    io_outs_101,
  output [5:0]    io_outs_100,
  output [5:0]    io_outs_99,
  output [5:0]    io_outs_98,
  output [5:0]    io_outs_97,
  output [5:0]    io_outs_96,
  output [5:0]    io_outs_95,
  output [5:0]    io_outs_94,
  output [5:0]    io_outs_93,
  output [5:0]    io_outs_92,
  output [5:0]    io_outs_91,
  output [5:0]    io_outs_90,
  output [5:0]    io_outs_89,
  output [5:0]    io_outs_88,
  output [5:0]    io_outs_87,
  output [5:0]    io_outs_86,
  output [5:0]    io_outs_85,
  output [5:0]    io_outs_84,
  output [5:0]    io_outs_83,
  output [5:0]    io_outs_82,
  output [5:0]    io_outs_81,
  output [5:0]    io_outs_80,
  output [5:0]    io_outs_79,
  output [5:0]    io_outs_78,
  output [5:0]    io_outs_77,
  output [5:0]    io_outs_76,
  output [5:0]    io_outs_75,
  output [5:0]    io_outs_74,
  output [5:0]    io_outs_73,
  output [5:0]    io_outs_72,
  output [5:0]    io_outs_71,
  output [5:0]    io_outs_70,
  output [5:0]    io_outs_69,
  output [5:0]    io_outs_68,
  output [5:0]    io_outs_67,
  output [5:0]    io_outs_66,
  output [5:0]    io_outs_65,
  output [5:0]    io_outs_64,
  output [5:0]    io_outs_63,
  output [5:0]    io_outs_62,
  output [5:0]    io_outs_61,
  output [5:0]    io_outs_60,
  output [5:0]    io_outs_59,
  output [5:0]    io_outs_58,
  output [5:0]    io_outs_57,
  output [5:0]    io_outs_56,
  output [5:0]    io_outs_55,
  output [5:0]    io_outs_54,
  output [5:0]    io_outs_53,
  output [5:0]    io_outs_52,
  output [5:0]    io_outs_51,
  output [5:0]    io_outs_50,
  output [5:0]    io_outs_49,
  output [5:0]    io_outs_48,
  output [5:0]    io_outs_47,
  output [5:0]    io_outs_46,
  output [5:0]    io_outs_45,
  output [5:0]    io_outs_44,
  output [5:0]    io_outs_43,
  output [5:0]    io_outs_42,
  output [5:0]    io_outs_41,
  output [5:0]    io_outs_40,
  output [5:0]    io_outs_39,
  output [5:0]    io_outs_38,
  output [5:0]    io_outs_37,
  output [5:0]    io_outs_36,
  output [5:0]    io_outs_35,
  output [5:0]    io_outs_34,
  output [5:0]    io_outs_33,
  output [5:0]    io_outs_32,
  output [5:0]    io_outs_31,
  output [5:0]    io_outs_30,
  output [5:0]    io_outs_29,
  output [5:0]    io_outs_28,
  output [5:0]    io_outs_27,
  output [5:0]    io_outs_26,
  output [5:0]    io_outs_25,
  output [5:0]    io_outs_24,
  output [5:0]    io_outs_23,
  output [5:0]    io_outs_22,
  output [5:0]    io_outs_21,
  output [5:0]    io_outs_20,
  output [5:0]    io_outs_19,
  output [5:0]    io_outs_18,
  output [5:0]    io_outs_17,
  output [5:0]    io_outs_16,
  output [5:0]    io_outs_15,
  output [5:0]    io_outs_14,
  output [5:0]    io_outs_13,
  output [5:0]    io_outs_12,
  output [5:0]    io_outs_11,
  output [5:0]    io_outs_10,
  output [5:0]    io_outs_9,
  output [5:0]    io_outs_8,
  output [5:0]    io_outs_7,
  output [5:0]    io_outs_6,
  output [5:0]    io_outs_5,
  output [5:0]    io_outs_4,
  output [5:0]    io_outs_3,
  output [5:0]    io_outs_2,
  output [5:0]    io_outs_1,
  output [5:0]    io_outs_0
);
  assign io_outs_191 = io_configuration[1151:1146]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_190 = io_configuration[1145:1140]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_189 = io_configuration[1139:1134]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_188 = io_configuration[1133:1128]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_187 = io_configuration[1127:1122]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_186 = io_configuration[1121:1116]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_185 = io_configuration[1115:1110]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_184 = io_configuration[1109:1104]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_183 = io_configuration[1103:1098]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_182 = io_configuration[1097:1092]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_181 = io_configuration[1091:1086]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_180 = io_configuration[1085:1080]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_179 = io_configuration[1079:1074]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_178 = io_configuration[1073:1068]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_177 = io_configuration[1067:1062]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_176 = io_configuration[1061:1056]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_175 = io_configuration[1055:1050]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_174 = io_configuration[1049:1044]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_173 = io_configuration[1043:1038]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_172 = io_configuration[1037:1032]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_171 = io_configuration[1031:1026]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_170 = io_configuration[1025:1020]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_169 = io_configuration[1019:1014]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_168 = io_configuration[1013:1008]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_167 = io_configuration[1007:1002]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_166 = io_configuration[1001:996]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_165 = io_configuration[995:990]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_164 = io_configuration[989:984]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_163 = io_configuration[983:978]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_162 = io_configuration[977:972]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_161 = io_configuration[971:966]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_160 = io_configuration[965:960]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_159 = io_configuration[959:954]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_158 = io_configuration[953:948]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_157 = io_configuration[947:942]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_156 = io_configuration[941:936]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_155 = io_configuration[935:930]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_154 = io_configuration[929:924]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_153 = io_configuration[923:918]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_152 = io_configuration[917:912]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_151 = io_configuration[911:906]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_150 = io_configuration[905:900]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_149 = io_configuration[899:894]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_148 = io_configuration[893:888]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_147 = io_configuration[887:882]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_146 = io_configuration[881:876]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_145 = io_configuration[875:870]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_144 = io_configuration[869:864]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_143 = io_configuration[863:858]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_142 = io_configuration[857:852]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_141 = io_configuration[851:846]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_140 = io_configuration[845:840]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_139 = io_configuration[839:834]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_138 = io_configuration[833:828]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_137 = io_configuration[827:822]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_136 = io_configuration[821:816]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_135 = io_configuration[815:810]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_134 = io_configuration[809:804]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_133 = io_configuration[803:798]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_132 = io_configuration[797:792]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_131 = io_configuration[791:786]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_130 = io_configuration[785:780]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_129 = io_configuration[779:774]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_128 = io_configuration[773:768]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_127 = io_configuration[767:762]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_126 = io_configuration[761:756]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_125 = io_configuration[755:750]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_124 = io_configuration[749:744]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_123 = io_configuration[743:738]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_122 = io_configuration[737:732]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_121 = io_configuration[731:726]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_120 = io_configuration[725:720]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_119 = io_configuration[719:714]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_118 = io_configuration[713:708]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_117 = io_configuration[707:702]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_116 = io_configuration[701:696]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_115 = io_configuration[695:690]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_114 = io_configuration[689:684]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_113 = io_configuration[683:678]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_112 = io_configuration[677:672]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_111 = io_configuration[671:666]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_110 = io_configuration[665:660]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_109 = io_configuration[659:654]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_108 = io_configuration[653:648]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_107 = io_configuration[647:642]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_106 = io_configuration[641:636]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_105 = io_configuration[635:630]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_104 = io_configuration[629:624]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_103 = io_configuration[623:618]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_102 = io_configuration[617:612]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_101 = io_configuration[611:606]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_100 = io_configuration[605:600]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_99 = io_configuration[599:594]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_98 = io_configuration[593:588]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_97 = io_configuration[587:582]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_96 = io_configuration[581:576]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_95 = io_configuration[575:570]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_94 = io_configuration[569:564]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_93 = io_configuration[563:558]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_92 = io_configuration[557:552]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_91 = io_configuration[551:546]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_90 = io_configuration[545:540]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_89 = io_configuration[539:534]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_88 = io_configuration[533:528]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_87 = io_configuration[527:522]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_86 = io_configuration[521:516]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_85 = io_configuration[515:510]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_84 = io_configuration[509:504]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_83 = io_configuration[503:498]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_82 = io_configuration[497:492]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_81 = io_configuration[491:486]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_80 = io_configuration[485:480]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_79 = io_configuration[479:474]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_78 = io_configuration[473:468]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_77 = io_configuration[467:462]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_76 = io_configuration[461:456]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_75 = io_configuration[455:450]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_74 = io_configuration[449:444]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_73 = io_configuration[443:438]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_72 = io_configuration[437:432]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_71 = io_configuration[431:426]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_70 = io_configuration[425:420]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_69 = io_configuration[419:414]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_68 = io_configuration[413:408]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_67 = io_configuration[407:402]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_66 = io_configuration[401:396]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_65 = io_configuration[395:390]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_64 = io_configuration[389:384]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_63 = io_configuration[383:378]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_62 = io_configuration[377:372]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_61 = io_configuration[371:366]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_60 = io_configuration[365:360]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_59 = io_configuration[359:354]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_58 = io_configuration[353:348]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_57 = io_configuration[347:342]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_56 = io_configuration[341:336]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_55 = io_configuration[335:330]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_54 = io_configuration[329:324]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_53 = io_configuration[323:318]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_52 = io_configuration[317:312]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_51 = io_configuration[311:306]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_50 = io_configuration[305:300]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_49 = io_configuration[299:294]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_48 = io_configuration[293:288]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_47 = io_configuration[287:282]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_46 = io_configuration[281:276]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_45 = io_configuration[275:270]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_44 = io_configuration[269:264]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_43 = io_configuration[263:258]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_42 = io_configuration[257:252]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_41 = io_configuration[251:246]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_40 = io_configuration[245:240]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_39 = io_configuration[239:234]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_38 = io_configuration[233:228]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_37 = io_configuration[227:222]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_36 = io_configuration[221:216]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_35 = io_configuration[215:210]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_34 = io_configuration[209:204]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_33 = io_configuration[203:198]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_32 = io_configuration[197:192]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_31 = io_configuration[191:186]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_30 = io_configuration[185:180]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_29 = io_configuration[179:174]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_28 = io_configuration[173:168]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_27 = io_configuration[167:162]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_26 = io_configuration[161:156]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_25 = io_configuration[155:150]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_24 = io_configuration[149:144]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_23 = io_configuration[143:138]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_22 = io_configuration[137:132]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_21 = io_configuration[131:126]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_20 = io_configuration[125:120]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_19 = io_configuration[119:114]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_18 = io_configuration[113:108]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_17 = io_configuration[107:102]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_16 = io_configuration[101:96]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_15 = io_configuration[95:90]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_14 = io_configuration[89:84]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_13 = io_configuration[83:78]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_12 = io_configuration[77:72]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_11 = io_configuration[71:66]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_10 = io_configuration[65:60]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_9 = io_configuration[59:54]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_8 = io_configuration[53:48]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_7 = io_configuration[47:42]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_6 = io_configuration[41:36]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_5 = io_configuration[35:30]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_4 = io_configuration[29:24]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_3 = io_configuration[23:18]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_2 = io_configuration[17:12]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_1 = io_configuration[11:6]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[5:0]; // @[BasicChiselModules.scala 490:18]
endmodule
module RegNextN(
  input         clock,
  input         reset,
  input  [2:0]  io_latency,
  input  [31:0] io_input,
  output [31:0] io_out
);
  reg [31:0] regArray_0; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_0;
  reg [31:0] regArray_1; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_1;
  reg [31:0] regArray_2; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_2;
  reg [31:0] regArray_3; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_3;
  reg [2:0] posReg; // @[BasicChiselModules.scala 41:23]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[BasicChiselModules.scala 43:19]
  wire [2:0] _T_3; // @[BasicChiselModules.scala 44:31]
  wire [1:0] _T_4;
  wire [31:0] _GEN_1; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_3; // @[BasicChiselModules.scala 44:12]
  wire [1:0] _T_5;
  wire [2:0] _T_7; // @[BasicChiselModules.scala 49:20]
  assign _T_1 = io_latency > 3'h0; // @[BasicChiselModules.scala 43:19]
  assign _T_3 = posReg - io_latency; // @[BasicChiselModules.scala 44:31]
  assign _T_4 = _T_3[1:0];
  assign _GEN_1 = 2'h1 == _T_4 ? regArray_1 : regArray_0; // @[BasicChiselModules.scala 44:12]
  assign _GEN_2 = 2'h2 == _T_4 ? regArray_2 : _GEN_1; // @[BasicChiselModules.scala 44:12]
  assign _GEN_3 = 2'h3 == _T_4 ? regArray_3 : _GEN_2; // @[BasicChiselModules.scala 44:12]
  assign _T_5 = posReg[1:0];
  assign _T_7 = posReg + 3'h1; // @[BasicChiselModules.scala 49:20]
  assign io_out = _T_1 ? _GEN_3 : io_input; // @[BasicChiselModules.scala 44:12 BasicChiselModules.scala 47:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regArray_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regArray_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regArray_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regArray_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  posReg = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regArray_0 <= 32'h0;
    end else if (_T_1) begin
      if (2'h0 == _T_5) begin
        regArray_0 <= io_input;
      end
    end
    if (reset) begin
      regArray_1 <= 32'h0;
    end else if (_T_1) begin
      if (2'h1 == _T_5) begin
        regArray_1 <= io_input;
      end
    end
    if (reset) begin
      regArray_2 <= 32'h0;
    end else if (_T_1) begin
      if (2'h2 == _T_5) begin
        regArray_2 <= io_input;
      end
    end
    if (reset) begin
      regArray_3 <= 32'h0;
    end else if (_T_1) begin
      if (2'h3 == _T_5) begin
        regArray_3 <= io_input;
      end
    end
    if (reset) begin
      posReg <= 3'h0;
    end else begin
      posReg <= _T_7;
    end
  end
endmodule
module Synchronizer(
  input         clock,
  input         reset,
  input  [3:0]  io_skewing,
  input  [31:0] io_input0,
  input  [31:0] io_input1,
  output [31:0] io_skewedInput0,
  output [31:0] io_skewedInput1
);
  wire  regNextN_clock; // @[BasicChiselModules.scala 66:24]
  wire  regNextN_reset; // @[BasicChiselModules.scala 66:24]
  wire [2:0] regNextN_io_latency; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_input; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_out; // @[BasicChiselModules.scala 66:24]
  wire  signal; // @[BasicChiselModules.scala 68:26]
  RegNextN regNextN ( // @[BasicChiselModules.scala 66:24]
    .clock(regNextN_clock),
    .reset(regNextN_reset),
    .io_latency(regNextN_io_latency),
    .io_input(regNextN_io_input),
    .io_out(regNextN_io_out)
  );
  assign signal = io_skewing[3]; // @[BasicChiselModules.scala 68:26]
  assign io_skewedInput0 = signal ? regNextN_io_out : io_input0; // @[BasicChiselModules.scala 73:21 BasicChiselModules.scala 78:21]
  assign io_skewedInput1 = signal ? io_input1 : regNextN_io_out; // @[BasicChiselModules.scala 74:21 BasicChiselModules.scala 77:21]
  assign regNextN_clock = clock;
  assign regNextN_reset = reset;
  assign regNextN_io_latency = io_skewing[2:0]; // @[BasicChiselModules.scala 69:23]
  assign regNextN_io_input = signal ? io_input0 : io_input1; // @[BasicChiselModules.scala 72:23 BasicChiselModules.scala 76:23]
endmodule
module Alu(
  input         clock,
  input         reset,
  input         io_en,
  input  [3:0]  io_skewing,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  Synchronizer_clock; // @[BasicChiselModules.scala 257:32]
  wire  Synchronizer_reset; // @[BasicChiselModules.scala 257:32]
  wire [3:0] Synchronizer_io_skewing; // @[BasicChiselModules.scala 257:32]
  wire [31:0] Synchronizer_io_input0; // @[BasicChiselModules.scala 257:32]
  wire [31:0] Synchronizer_io_input1; // @[BasicChiselModules.scala 257:32]
  wire [31:0] Synchronizer_io_skewedInput0; // @[BasicChiselModules.scala 257:32]
  wire [31:0] Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 257:32]
  wire [31:0] _T_1; // @[BasicChiselModules.scala 230:55]
  wire [31:0] _T_3; // @[BasicChiselModules.scala 231:55]
  wire [31:0] _T_4; // @[BasicChiselModules.scala 232:55]
  wire [31:0] _T_5; // @[BasicChiselModules.scala 233:54]
  wire [31:0] _T_6; // @[BasicChiselModules.scala 234:55]
  wire [63:0] _T_7; // @[BasicChiselModules.scala 235:55]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [63:0] _T_13; // @[Mux.scala 68:16]
  wire  _T_14; // @[Mux.scala 68:19]
  wire [63:0] _T_15; // @[Mux.scala 68:16]
  wire  _T_16; // @[Mux.scala 68:19]
  wire [63:0] _T_17; // @[Mux.scala 68:16]
  wire  _T_18; // @[Mux.scala 68:19]
  wire [63:0] _T_19; // @[Mux.scala 68:16]
  wire  _T_20; // @[Mux.scala 68:19]
  wire [63:0] _T_21; // @[Mux.scala 68:16]
  wire  _T_22; // @[Mux.scala 68:19]
  wire [63:0] _T_23; // @[Mux.scala 68:16]
  wire [63:0] _GEN_0; // @[BasicChiselModules.scala 283:15]
  Synchronizer Synchronizer ( // @[BasicChiselModules.scala 257:32]
    .clock(Synchronizer_clock),
    .reset(Synchronizer_reset),
    .io_skewing(Synchronizer_io_skewing),
    .io_input0(Synchronizer_io_input0),
    .io_input1(Synchronizer_io_input1),
    .io_skewedInput0(Synchronizer_io_skewedInput0),
    .io_skewedInput1(Synchronizer_io_skewedInput1)
  );
  assign _T_1 = Synchronizer_io_skewedInput0 + Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 230:55]
  assign _T_3 = Synchronizer_io_skewedInput0 - Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 231:55]
  assign _T_4 = Synchronizer_io_skewedInput0 & Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 232:55]
  assign _T_5 = Synchronizer_io_skewedInput0 | Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 233:54]
  assign _T_6 = Synchronizer_io_skewedInput0 ^ Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 234:55]
  assign _T_7 = Synchronizer_io_skewedInput0 * Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 235:55]
  assign _T_9 = Synchronizer_io_skewedInput1; // @[Mux.scala 68:16]
  assign _T_10 = 4'hc == io_configuration; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? Synchronizer_io_skewedInput0 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 4'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_13 = _T_12 ? _T_7 : {{32'd0}, _T_11}; // @[Mux.scala 68:16]
  assign _T_14 = 4'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_15 = _T_14 ? {{32'd0}, _T_6} : _T_13; // @[Mux.scala 68:16]
  assign _T_16 = 4'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_17 = _T_16 ? {{32'd0}, _T_5} : _T_15; // @[Mux.scala 68:16]
  assign _T_18 = 4'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_19 = _T_18 ? {{32'd0}, _T_4} : _T_17; // @[Mux.scala 68:16]
  assign _T_20 = 4'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_21 = _T_20 ? {{32'd0}, _T_3} : _T_19; // @[Mux.scala 68:16]
  assign _T_22 = 4'h0 == io_configuration; // @[Mux.scala 68:19]
  assign _T_23 = _T_22 ? {{32'd0}, _T_1} : _T_21; // @[Mux.scala 68:16]
  assign _GEN_0 = io_en ? _T_23 : 64'h0; // @[BasicChiselModules.scala 283:15]
  assign io_outs_0 = _GEN_0[31:0]; // @[BasicChiselModules.scala 284:9 BasicChiselModules.scala 287:11]
  assign Synchronizer_clock = clock;
  assign Synchronizer_reset = reset;
  assign Synchronizer_io_skewing = io_skewing; // @[BasicChiselModules.scala 261:31]
  assign Synchronizer_io_input0 = io_inputs_0; // @[BasicChiselModules.scala 258:30]
  assign Synchronizer_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 259:30]
endmodule
module ScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [1:0] io_waitCycle,
  output       io_valid
);
  reg  state; // @[BasicChiselModules.scala 139:22]
  reg [31:0] _RAND_0;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 140:21]
  reg [31:0] _RAND_1;
  wire  _T; // @[BasicChiselModules.scala 142:25]
  wire  _T_2; // @[BasicChiselModules.scala 145:16]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 149:30]
  wire  _GEN_0; // @[BasicChiselModules.scala 146:39]
  wire  _GEN_2; // @[BasicChiselModules.scala 145:28]
  wire  _GEN_4; // @[BasicChiselModules.scala 144:15]
  assign _T = cycleReg == io_waitCycle; // @[BasicChiselModules.scala 142:25]
  assign _T_2 = state == 1'h0; // @[BasicChiselModules.scala 145:16]
  assign _T_5 = cycleReg + 2'h1; // @[BasicChiselModules.scala 149:30]
  assign _GEN_0 = _T | state; // @[BasicChiselModules.scala 146:39]
  assign _GEN_2 = _T_2 ? _GEN_0 : state; // @[BasicChiselModules.scala 145:28]
  assign _GEN_4 = io_en & _GEN_2; // @[BasicChiselModules.scala 144:15]
  assign io_valid = _T & io_en; // @[BasicChiselModules.scala 142:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_4;
    end
    if (io_en) begin
      if (_T_2) begin
        if (!(_T)) begin
          cycleReg <= _T_5;
        end
      end
    end else begin
      cycleReg <= 2'h0;
    end
  end
endmodule
module MultiIIScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [5:0] io_schedules_0,
  input  [5:0] io_schedules_1,
  input  [5:0] io_schedules_2,
  input  [5:0] io_schedules_3,
  input  [5:0] io_schedules_4,
  input  [5:0] io_schedules_5,
  input  [5:0] io_schedules_6,
  input  [5:0] io_schedules_7,
  input  [2:0] io_II,
  output       io_valid,
  output [3:0] io_skewing
);
  wire  ScheduleController_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_1_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_1_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_1_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_1_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_1_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_2_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_2_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_2_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_2_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_2_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_3_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_3_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_3_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_3_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_3_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_4_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_4_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_4_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_4_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_4_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_5_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_5_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_5_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_5_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_5_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_6_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_6_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_6_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_6_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_6_io_valid; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_7_clock; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_7_reset; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_7_io_en; // @[BasicChiselModules.scala 174:79]
  wire [1:0] ScheduleController_7_io_waitCycle; // @[BasicChiselModules.scala 174:79]
  wire  ScheduleController_7_io_valid; // @[BasicChiselModules.scala 174:79]
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 171:25]
  reg [31:0] _RAND_0;
  reg  _T_1_0; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_1;
  reg  _T_1_1; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_2;
  reg  _T_1_2; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_3;
  reg  _T_1_3; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_4;
  reg  _T_1_4; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_5;
  reg  _T_1_5; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_6;
  reg  _T_1_6; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_7;
  reg  _T_1_7; // @[BasicChiselModules.scala 175:28]
  reg [31:0] _RAND_8;
  wire  _GEN_1; // @[BasicChiselModules.scala 182:14]
  wire  _GEN_2; // @[BasicChiselModules.scala 182:14]
  wire  _GEN_3; // @[BasicChiselModules.scala 182:14]
  wire  _GEN_4; // @[BasicChiselModules.scala 182:14]
  wire  _GEN_5; // @[BasicChiselModules.scala 182:14]
  wire  _GEN_6; // @[BasicChiselModules.scala 182:14]
  wire [5:0] _GEN_9; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_10; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_11; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_12; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_13; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_14; // @[BasicChiselModules.scala 189:41]
  wire [5:0] _GEN_15; // @[BasicChiselModules.scala 189:41]
  wire [2:0] _T_13; // @[BasicChiselModules.scala 195:29]
  wire  _T_14; // @[BasicChiselModules.scala 195:19]
  wire [2:0] _T_16; // @[BasicChiselModules.scala 198:28]
  ScheduleController ScheduleController ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_clock),
    .reset(ScheduleController_reset),
    .io_en(ScheduleController_io_en),
    .io_waitCycle(ScheduleController_io_waitCycle),
    .io_valid(ScheduleController_io_valid)
  );
  ScheduleController ScheduleController_1 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_1_clock),
    .reset(ScheduleController_1_reset),
    .io_en(ScheduleController_1_io_en),
    .io_waitCycle(ScheduleController_1_io_waitCycle),
    .io_valid(ScheduleController_1_io_valid)
  );
  ScheduleController ScheduleController_2 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_2_clock),
    .reset(ScheduleController_2_reset),
    .io_en(ScheduleController_2_io_en),
    .io_waitCycle(ScheduleController_2_io_waitCycle),
    .io_valid(ScheduleController_2_io_valid)
  );
  ScheduleController ScheduleController_3 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_3_clock),
    .reset(ScheduleController_3_reset),
    .io_en(ScheduleController_3_io_en),
    .io_waitCycle(ScheduleController_3_io_waitCycle),
    .io_valid(ScheduleController_3_io_valid)
  );
  ScheduleController ScheduleController_4 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_4_clock),
    .reset(ScheduleController_4_reset),
    .io_en(ScheduleController_4_io_en),
    .io_waitCycle(ScheduleController_4_io_waitCycle),
    .io_valid(ScheduleController_4_io_valid)
  );
  ScheduleController ScheduleController_5 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_5_clock),
    .reset(ScheduleController_5_reset),
    .io_en(ScheduleController_5_io_en),
    .io_waitCycle(ScheduleController_5_io_waitCycle),
    .io_valid(ScheduleController_5_io_valid)
  );
  ScheduleController ScheduleController_6 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_6_clock),
    .reset(ScheduleController_6_reset),
    .io_en(ScheduleController_6_io_en),
    .io_waitCycle(ScheduleController_6_io_waitCycle),
    .io_valid(ScheduleController_6_io_valid)
  );
  ScheduleController ScheduleController_7 ( // @[BasicChiselModules.scala 174:79]
    .clock(ScheduleController_7_clock),
    .reset(ScheduleController_7_reset),
    .io_en(ScheduleController_7_io_en),
    .io_waitCycle(ScheduleController_7_io_waitCycle),
    .io_valid(ScheduleController_7_io_valid)
  );
  assign _GEN_1 = 3'h1 == cycleReg ? _T_1_1 : _T_1_0; // @[BasicChiselModules.scala 182:14]
  assign _GEN_2 = 3'h2 == cycleReg ? _T_1_2 : _GEN_1; // @[BasicChiselModules.scala 182:14]
  assign _GEN_3 = 3'h3 == cycleReg ? _T_1_3 : _GEN_2; // @[BasicChiselModules.scala 182:14]
  assign _GEN_4 = 3'h4 == cycleReg ? _T_1_4 : _GEN_3; // @[BasicChiselModules.scala 182:14]
  assign _GEN_5 = 3'h5 == cycleReg ? _T_1_5 : _GEN_4; // @[BasicChiselModules.scala 182:14]
  assign _GEN_6 = 3'h6 == cycleReg ? _T_1_6 : _GEN_5; // @[BasicChiselModules.scala 182:14]
  assign _GEN_9 = 3'h1 == cycleReg ? io_schedules_1 : io_schedules_0; // @[BasicChiselModules.scala 189:41]
  assign _GEN_10 = 3'h2 == cycleReg ? io_schedules_2 : _GEN_9; // @[BasicChiselModules.scala 189:41]
  assign _GEN_11 = 3'h3 == cycleReg ? io_schedules_3 : _GEN_10; // @[BasicChiselModules.scala 189:41]
  assign _GEN_12 = 3'h4 == cycleReg ? io_schedules_4 : _GEN_11; // @[BasicChiselModules.scala 189:41]
  assign _GEN_13 = 3'h5 == cycleReg ? io_schedules_5 : _GEN_12; // @[BasicChiselModules.scala 189:41]
  assign _GEN_14 = 3'h6 == cycleReg ? io_schedules_6 : _GEN_13; // @[BasicChiselModules.scala 189:41]
  assign _GEN_15 = 3'h7 == cycleReg ? io_schedules_7 : _GEN_14; // @[BasicChiselModules.scala 189:41]
  assign _T_13 = io_II - 3'h1; // @[BasicChiselModules.scala 195:29]
  assign _T_14 = cycleReg == _T_13; // @[BasicChiselModules.scala 195:19]
  assign _T_16 = cycleReg + 3'h1; // @[BasicChiselModules.scala 198:28]
  assign io_valid = 3'h7 == cycleReg ? _T_1_7 : _GEN_6; // @[BasicChiselModules.scala 182:14]
  assign io_skewing = _GEN_15[5:2]; // @[BasicChiselModules.scala 189:16]
  assign ScheduleController_clock = clock;
  assign ScheduleController_reset = reset;
  assign ScheduleController_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_io_waitCycle = io_schedules_0[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_1_clock = clock;
  assign ScheduleController_1_reset = reset;
  assign ScheduleController_1_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_1_io_waitCycle = io_schedules_1[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_2_clock = clock;
  assign ScheduleController_2_reset = reset;
  assign ScheduleController_2_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_2_io_waitCycle = io_schedules_2[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_3_clock = clock;
  assign ScheduleController_3_reset = reset;
  assign ScheduleController_3_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_3_io_waitCycle = io_schedules_3[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_4_clock = clock;
  assign ScheduleController_4_reset = reset;
  assign ScheduleController_4_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_4_io_waitCycle = io_schedules_4[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_5_clock = clock;
  assign ScheduleController_5_reset = reset;
  assign ScheduleController_5_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_5_io_waitCycle = io_schedules_5[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_6_clock = clock;
  assign ScheduleController_6_reset = reset;
  assign ScheduleController_6_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_6_io_waitCycle = io_schedules_6[1:0]; // @[BasicChiselModules.scala 179:39]
  assign ScheduleController_7_clock = clock;
  assign ScheduleController_7_reset = reset;
  assign ScheduleController_7_io_en = io_en; // @[BasicChiselModules.scala 178:32]
  assign ScheduleController_7_io_waitCycle = io_schedules_7[1:0]; // @[BasicChiselModules.scala 179:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleReg = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1_3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1_4 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1_6 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1_7 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleReg <= 3'h7;
    end else if (io_en) begin
      if (_T_14) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_16;
      end
    end
    if (reset) begin
      _T_1_0 <= 1'h0;
    end else begin
      _T_1_0 <= ScheduleController_io_valid;
    end
    if (reset) begin
      _T_1_1 <= 1'h0;
    end else begin
      _T_1_1 <= ScheduleController_1_io_valid;
    end
    if (reset) begin
      _T_1_2 <= 1'h0;
    end else begin
      _T_1_2 <= ScheduleController_2_io_valid;
    end
    if (reset) begin
      _T_1_3 <= 1'h0;
    end else begin
      _T_1_3 <= ScheduleController_3_io_valid;
    end
    if (reset) begin
      _T_1_4 <= 1'h0;
    end else begin
      _T_1_4 <= ScheduleController_4_io_valid;
    end
    if (reset) begin
      _T_1_5 <= 1'h0;
    end else begin
      _T_1_5 <= ScheduleController_5_io_valid;
    end
    if (reset) begin
      _T_1_6 <= 1'h0;
    end else begin
      _T_1_6 <= ScheduleController_6_io_valid;
    end
    if (reset) begin
      _T_1_7 <= 1'h0;
    end else begin
      _T_1_7 <= ScheduleController_7_io_valid;
    end
  end
endmodule
module Dispatch_1(
  input  [1:0] io_configuration,
  output       io_outs_1,
  output       io_outs_0
);
  assign io_outs_1 = io_configuration[1]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[0]; // @[BasicChiselModules.scala 490:18]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire [1:0] Dispatch_io_configuration; // @[BasicChiselModules.scala 358:26]
  wire  Dispatch_io_outs_1; // @[BasicChiselModules.scala 358:26]
  wire  Dispatch_io_outs_0; // @[BasicChiselModules.scala 358:26]
  wire  _T_1; // @[BasicChiselModules.scala 362:37]
  reg [31:0] _T_3_0; // @[BasicChiselModules.scala 364:23]
  reg [31:0] _RAND_0;
  reg [31:0] _T_3_1; // @[BasicChiselModules.scala 364:23]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[BasicChiselModules.scala 366:20]
  Dispatch_1 Dispatch ( // @[BasicChiselModules.scala 358:26]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  assign _T_1 = io_configuration[2]; // @[BasicChiselModules.scala 362:37]
  assign _T_4 = _T_1 == 1'h0; // @[BasicChiselModules.scala 366:20]
  assign io_outs_0 = Dispatch_io_outs_1 ? _T_3_1 : _T_3_0; // @[BasicChiselModules.scala 372:18]
  assign Dispatch_io_configuration = io_configuration[1:0]; // @[BasicChiselModules.scala 360:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3_0 <= 32'h0;
    end else if (_T_4) begin
      if (1'h0 == Dispatch_io_outs_0) begin
        _T_3_0 <= io_inputs_0;
      end
    end
    if (reset) begin
      _T_3_1 <= 32'h0;
    end else if (_T_4) begin
      if (Dispatch_io_outs_0) begin
        _T_3_1 <= io_inputs_0;
      end
    end
  end
endmodule
module Multiplexer(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  assign _T = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_4 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_3 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_1 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_8 ? io_inputs_0 : _T_7; // @[BasicChiselModules.scala 396:14]
endmodule
module Multiplexer_5(
  input         io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  assign _T_1 = io_configuration ? io_inputs_1 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 1'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_2 ? io_inputs_0 : _T_1; // @[BasicChiselModules.scala 396:14]
endmodule
module Multiplexer_8(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  assign _T = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_5 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_4 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_3 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_2 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_1 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_10 ? io_inputs_0 : _T_9; // @[BasicChiselModules.scala 396:14]
endmodule
module ConstUnit(
  input  [31:0] io_configuration,
  output [31:0] io_outs_0
);
  assign io_outs_0 = io_configuration; // @[BasicChiselModules.scala 429:14]
endmodule
module SimpleDualPortSram(
  input         clock,
  input         io_a_en,
  input         io_a_we,
  input  [5:0]  io_a_addr,
  input  [31:0] io_a_din,
  input         io_b_en,
  input  [5:0]  io_b_addr,
  output [31:0] io_b_dout
);
  reg [31:0] mem [0:63]; // @[Mem.scala 201:16]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_2_data; // @[Mem.scala 201:16]
  wire [5:0] mem__T_2_addr; // @[Mem.scala 201:16]
  wire [31:0] mem__T_1_data; // @[Mem.scala 201:16]
  wire [5:0] mem__T_1_addr; // @[Mem.scala 201:16]
  wire  mem__T_1_mask; // @[Mem.scala 201:16]
  wire  mem__T_1_en; // @[Mem.scala 201:16]
  reg [31:0] dout; // @[Mem.scala 202:17]
  reg [31:0] _RAND_1;
  assign mem__T_2_addr = io_b_addr;
  assign mem__T_2_data = mem[mem__T_2_addr]; // @[Mem.scala 201:16]
  assign mem__T_1_data = io_a_din;
  assign mem__T_1_addr = io_a_addr;
  assign mem__T_1_mask = 1'h1;
  assign mem__T_1_en = io_a_en & io_a_we;
  assign io_b_dout = dout; // @[Mem.scala 204:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dout = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_1_en & mem__T_1_mask) begin
      mem[mem__T_1_addr] <= mem__T_1_data; // @[Mem.scala 201:16]
    end
    if (io_b_en) begin
      dout <= mem__T_2_data;
    end
  end
endmodule
module EnqMem(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_mem_en,
  output        io_mem_we,
  output [5:0]  io_mem_addr,
  output [31:0] io_mem_din,
  input  [5:0]  io_base,
  input         io_en,
  input         io_start,
  output        io_idle
);
  reg  state; // @[EnqMem.scala 64:22]
  reg [31:0] _RAND_0;
  reg [5:0] mem_index; // @[EnqMem.scala 68:22]
  reg [31:0] _RAND_1;
  reg [31:0] data_in; // @[EnqMem.scala 69:20]
  reg [31:0] _RAND_2;
  wire  _T; // @[EnqMem.scala 75:21]
  wire  _T_1; // @[EnqMem.scala 75:38]
  wire  _T_3; // @[EnqMem.scala 79:19]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire [5:0] _T_8; // @[EnqMem.scala 95:34]
  wire  _GEN_12; // @[EnqMem.scala 91:33]
  assign _T = state == 1'h0; // @[EnqMem.scala 75:21]
  assign _T_1 = io_in_valid == 1'h0; // @[EnqMem.scala 75:38]
  assign _T_3 = io_idle & io_start; // @[EnqMem.scala 79:19]
  assign _T_5 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = mem_index + 6'h1; // @[EnqMem.scala 95:34]
  assign _GEN_12 = state | _T; // @[EnqMem.scala 91:33]
  assign io_in_ready = io_en & _GEN_12; // @[Decoupled.scala 72:20 Decoupled.scala 65:20 Decoupled.scala 65:20]
  assign io_mem_en = io_en & state; // @[Mem.scala 73:8 Mem.scala 69:8]
  assign io_mem_we = io_en & state; // @[Mem.scala 74:8 Mem.scala 70:8]
  assign io_mem_addr = mem_index; // @[EnqMem.scala 93:23]
  assign io_mem_din = data_in; // @[EnqMem.scala 94:22]
  assign io_idle = _T & _T_1; // @[EnqMem.scala 75:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_index = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_in = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else if (io_en) begin
      if (state) begin
        state <= _T_5;
      end else if (_T) begin
        state <= _T_5;
      end else if (_T_3) begin
        state <= 1'h0;
      end
    end
    if (io_en) begin
      if (state) begin
        mem_index <= _T_8;
      end else if (_T_3) begin
        mem_index <= io_base;
      end
    end
    if (io_en) begin
      if (state) begin
        data_in <= io_in_bits;
      end else if (_T) begin
        data_in <= io_in_bits;
      end
    end
  end
endmodule
module Handshake(
  output       io_enq_ready,
  input        io_enq_valid,
  input  [5:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [5:0] io_deq_bits
);
  assign io_enq_ready = io_deq_ready; // @[BusHelper.scala 11:10]
  assign io_deq_valid = io_enq_valid; // @[BusHelper.scala 11:10]
  assign io_deq_bits = io_enq_bits; // @[BusHelper.scala 11:10]
endmodule
module Handshake_1(
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
  assign io_enq_ready = io_deq_ready; // @[BusHelper.scala 11:10]
  assign io_deq_valid = io_enq_valid; // @[BusHelper.scala 11:10]
  assign io_deq_bits = io_enq_bits; // @[BusHelper.scala 11:10]
endmodule
module EnqAddrDeqMem(
  input         clock,
  input         reset,
  output        io_iaddr_ready,
  input         io_iaddr_valid,
  input  [5:0]  io_iaddr_bits,
  output        io_mem_en,
  output [5:0]  io_mem_addr,
  input  [31:0] io_mem_dout,
  input         io_odata_ready,
  output        io_odata_valid,
  output [31:0] io_odata_bits,
  output        io_idle
);
  reg  token; // @[DeqMem.scala 216:22]
  reg [31:0] _RAND_0;
  wire  _T; // @[DeqMem.scala 223:21]
  wire  _T_1; // @[DeqMem.scala 223:53]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_0; // @[DeqMem.scala 232:27]
  wire  _GEN_4; // @[DeqMem.scala 230:15]
  wire  _T_4; // @[DeqMem.scala 238:19]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[DeqMem.scala 240:27]
  assign _T = token == 1'h0; // @[DeqMem.scala 223:21]
  assign _T_1 = io_iaddr_valid == 1'h0; // @[DeqMem.scala 223:53]
  assign _T_3 = io_odata_ready & io_odata_valid; // @[Decoupled.scala 40:37]
  assign _GEN_0 = _T_3 ? 1'h0 : token; // @[DeqMem.scala 232:27]
  assign _GEN_4 = token ? _GEN_0 : token; // @[DeqMem.scala 230:15]
  assign _T_4 = _GEN_4 == 1'h0; // @[DeqMem.scala 238:19]
  assign _T_5 = io_iaddr_ready & io_iaddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_5 | _GEN_4; // @[DeqMem.scala 240:27]
  assign io_iaddr_ready = _GEN_4 == 1'h0; // @[Decoupled.scala 72:20 Decoupled.scala 65:20]
  assign io_mem_en = _T_4 & _T_5; // @[Mem.scala 43:8 Mem.scala 40:8]
  assign io_mem_addr = io_iaddr_bits; // @[DeqMem.scala 243:19]
  assign io_odata_valid = token; // @[Decoupled.scala 56:20 Decoupled.scala 47:20]
  assign io_odata_bits = io_mem_dout; // @[Decoupled.scala 48:19]
  assign io_idle = _T & _T_1; // @[DeqMem.scala 223:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  token = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      token <= 1'h0;
    end else if (_T_4) begin
      token <= _GEN_6;
    end else if (token) begin
      if (_T_3) begin
        token <= 1'h0;
      end
    end
  end
endmodule
module DeqMem(
  input         clock,
  input         reset,
  output        io_mem_en,
  output [5:0]  io_mem_addr,
  input  [31:0] io_mem_dout,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits,
  input  [5:0]  io_base,
  input  [5:0]  io_len,
  input         io_en,
  input         io_start,
  output        io_idle
);
  wire  iaddr_hs_io_enq_ready; // @[DeqMem.scala 103:24]
  wire  iaddr_hs_io_enq_valid; // @[DeqMem.scala 103:24]
  wire [5:0] iaddr_hs_io_enq_bits; // @[DeqMem.scala 103:24]
  wire  iaddr_hs_io_deq_ready; // @[DeqMem.scala 103:24]
  wire  iaddr_hs_io_deq_valid; // @[DeqMem.scala 103:24]
  wire [5:0] iaddr_hs_io_deq_bits; // @[DeqMem.scala 103:24]
  wire  odata_hs_io_enq_ready; // @[DeqMem.scala 107:24]
  wire  odata_hs_io_enq_valid; // @[DeqMem.scala 107:24]
  wire [31:0] odata_hs_io_enq_bits; // @[DeqMem.scala 107:24]
  wire  odata_hs_io_deq_ready; // @[DeqMem.scala 107:24]
  wire  odata_hs_io_deq_valid; // @[DeqMem.scala 107:24]
  wire [31:0] odata_hs_io_deq_bits; // @[DeqMem.scala 107:24]
  wire  EnqAddrDeqMem_clock; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_reset; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_iaddr_ready; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_iaddr_valid; // @[DeqMem.scala 57:22]
  wire [5:0] EnqAddrDeqMem_io_iaddr_bits; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_mem_en; // @[DeqMem.scala 57:22]
  wire [5:0] EnqAddrDeqMem_io_mem_addr; // @[DeqMem.scala 57:22]
  wire [31:0] EnqAddrDeqMem_io_mem_dout; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_odata_ready; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_odata_valid; // @[DeqMem.scala 57:22]
  wire [31:0] EnqAddrDeqMem_io_odata_bits; // @[DeqMem.scala 57:22]
  wire  EnqAddrDeqMem_io_idle; // @[DeqMem.scala 57:22]
  reg [1:0] state; // @[DeqMem.scala 94:22]
  reg [31:0] _RAND_0;
  reg [5:0] mem_index; // @[DeqMem.scala 98:22]
  reg [31:0] _RAND_1;
  reg [31:0] mem_data; // @[DeqMem.scala 99:21]
  reg [31:0] _RAND_2;
  reg [5:0] remain; // @[DeqMem.scala 101:19]
  reg [31:0] _RAND_3;
  wire  _T_1; // @[DeqMem.scala 126:18]
  wire [5:0] _GEN_1; // @[DeqMem.scala 126:31]
  wire [5:0] _GEN_3; // @[DeqMem.scala 126:31]
  wire  _T_2; // @[DeqMem.scala 133:16]
  wire  _T_3; // @[DeqMem.scala 189:17]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire [5:0] _T_6; // @[DeqMem.scala 192:32]
  wire [5:0] _T_8; // @[DeqMem.scala 193:26]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[DeqMem.scala 200:27]
  wire  _GEN_12; // @[DeqMem.scala 133:29]
  wire  _T_11; // @[DeqMem.scala 139:20]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[DeqMem.scala 189:24]
  wire  _GEN_27; // @[DeqMem.scala 141:31]
  wire  _GEN_31; // @[DeqMem.scala 141:31]
  wire  _GEN_36; // @[DeqMem.scala 139:32]
  wire  _GEN_40; // @[DeqMem.scala 139:32]
  Handshake iaddr_hs ( // @[DeqMem.scala 103:24]
    .io_enq_ready(iaddr_hs_io_enq_ready),
    .io_enq_valid(iaddr_hs_io_enq_valid),
    .io_enq_bits(iaddr_hs_io_enq_bits),
    .io_deq_ready(iaddr_hs_io_deq_ready),
    .io_deq_valid(iaddr_hs_io_deq_valid),
    .io_deq_bits(iaddr_hs_io_deq_bits)
  );
  Handshake_1 odata_hs ( // @[DeqMem.scala 107:24]
    .io_enq_ready(odata_hs_io_enq_ready),
    .io_enq_valid(odata_hs_io_enq_valid),
    .io_enq_bits(odata_hs_io_enq_bits),
    .io_deq_ready(odata_hs_io_deq_ready),
    .io_deq_valid(odata_hs_io_deq_valid),
    .io_deq_bits(odata_hs_io_deq_bits)
  );
  EnqAddrDeqMem EnqAddrDeqMem ( // @[DeqMem.scala 57:22]
    .clock(EnqAddrDeqMem_clock),
    .reset(EnqAddrDeqMem_reset),
    .io_iaddr_ready(EnqAddrDeqMem_io_iaddr_ready),
    .io_iaddr_valid(EnqAddrDeqMem_io_iaddr_valid),
    .io_iaddr_bits(EnqAddrDeqMem_io_iaddr_bits),
    .io_mem_en(EnqAddrDeqMem_io_mem_en),
    .io_mem_addr(EnqAddrDeqMem_io_mem_addr),
    .io_mem_dout(EnqAddrDeqMem_io_mem_dout),
    .io_odata_ready(EnqAddrDeqMem_io_odata_ready),
    .io_odata_valid(EnqAddrDeqMem_io_odata_valid),
    .io_odata_bits(EnqAddrDeqMem_io_odata_bits),
    .io_idle(EnqAddrDeqMem_io_idle)
  );
  assign _T_1 = io_idle & io_start; // @[DeqMem.scala 126:18]
  assign _GEN_1 = _T_1 ? io_base : mem_index; // @[DeqMem.scala 126:31]
  assign _GEN_3 = _T_1 ? io_len : remain; // @[DeqMem.scala 126:31]
  assign _T_2 = state == 2'h1; // @[DeqMem.scala 133:16]
  assign _T_3 = remain > 6'h0; // @[DeqMem.scala 189:17]
  assign _T_4 = iaddr_hs_io_enq_ready & iaddr_hs_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = mem_index + 6'h1; // @[DeqMem.scala 192:32]
  assign _T_8 = remain - 6'h1; // @[DeqMem.scala 193:26]
  assign _T_9 = odata_hs_io_deq_ready & odata_hs_io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = EnqAddrDeqMem_io_idle == 1'h0; // @[DeqMem.scala 200:27]
  assign _GEN_12 = _T_2 & _T_3; // @[DeqMem.scala 133:29]
  assign _T_11 = state == 2'h2; // @[DeqMem.scala 139:20]
  assign _T_12 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_3 | _GEN_12; // @[DeqMem.scala 189:24]
  assign _GEN_27 = _T_12 ? _GEN_21 : _GEN_12; // @[DeqMem.scala 141:31]
  assign _GEN_31 = _T_12 | _T_2; // @[DeqMem.scala 141:31]
  assign _GEN_36 = _T_11 ? _GEN_27 : _GEN_12; // @[DeqMem.scala 139:32]
  assign _GEN_40 = _T_11 ? _GEN_31 : _T_2; // @[DeqMem.scala 139:32]
  assign io_mem_en = EnqAddrDeqMem_io_mem_en; // @[Mem.scala 43:8 DeqMem.scala 71:22]
  assign io_mem_addr = EnqAddrDeqMem_io_mem_addr; // @[DeqMem.scala 72:24]
  assign io_out_valid = io_en & _T_11; // @[Decoupled.scala 56:20 Decoupled.scala 47:20]
  assign io_out_bits = mem_data; // @[Decoupled.scala 48:19]
  assign io_idle = state == 2'h0; // @[DeqMem.scala 120:11]
  assign iaddr_hs_io_enq_valid = io_en & _GEN_36; // @[Decoupled.scala 56:20 Decoupled.scala 47:20 Decoupled.scala 47:20]
  assign iaddr_hs_io_enq_bits = mem_index; // @[Decoupled.scala 48:19 Decoupled.scala 48:19]
  assign iaddr_hs_io_deq_ready = EnqAddrDeqMem_io_iaddr_ready; // @[Decoupled.scala 72:20 DeqMem.scala 70:21]
  assign odata_hs_io_enq_valid = EnqAddrDeqMem_io_odata_valid; // @[Decoupled.scala 56:20 DeqMem.scala 74:21]
  assign odata_hs_io_enq_bits = EnqAddrDeqMem_io_odata_bits; // @[DeqMem.scala 74:21]
  assign odata_hs_io_deq_ready = io_en & _GEN_40; // @[Decoupled.scala 72:20 Decoupled.scala 65:20 Decoupled.scala 65:20]
  assign EnqAddrDeqMem_clock = clock;
  assign EnqAddrDeqMem_reset = reset;
  assign EnqAddrDeqMem_io_iaddr_valid = iaddr_hs_io_deq_valid; // @[Decoupled.scala 56:20 DeqMem.scala 70:21]
  assign EnqAddrDeqMem_io_iaddr_bits = iaddr_hs_io_deq_bits; // @[DeqMem.scala 70:21]
  assign EnqAddrDeqMem_io_mem_dout = io_mem_dout; // @[DeqMem.scala 73:24]
  assign EnqAddrDeqMem_io_odata_ready = odata_hs_io_enq_ready; // @[Decoupled.scala 72:20 DeqMem.scala 74:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_index = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  remain = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_9) begin
            state <= 2'h2;
          end else if (_T_10) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end else if (_T_2) begin
          if (_T_9) begin
            state <= 2'h2;
          end else if (_T_10) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end else if (_T_1) begin
          state <= 2'h1;
        end
      end else if (_T_2) begin
        if (_T_9) begin
          state <= 2'h2;
        end else if (_T_10) begin
          state <= 2'h1;
        end else begin
          state <= 2'h0;
        end
      end else if (_T_1) begin
        state <= 2'h1;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_3) begin
            if (_T_4) begin
              mem_index <= _T_6;
            end else if (_T_2) begin
              if (_T_3) begin
                if (_T_4) begin
                  mem_index <= _T_6;
                end else if (_T_1) begin
                  mem_index <= io_base;
                end
              end else if (_T_1) begin
                mem_index <= io_base;
              end
            end else if (_T_1) begin
              mem_index <= io_base;
            end
          end else if (_T_2) begin
            if (_T_3) begin
              if (_T_4) begin
                mem_index <= _T_6;
              end else if (_T_1) begin
                mem_index <= io_base;
              end
            end else begin
              mem_index <= _GEN_1;
            end
          end else begin
            mem_index <= _GEN_1;
          end
        end else if (_T_2) begin
          if (_T_3) begin
            if (_T_4) begin
              mem_index <= _T_6;
            end else begin
              mem_index <= _GEN_1;
            end
          end else begin
            mem_index <= _GEN_1;
          end
        end else begin
          mem_index <= _GEN_1;
        end
      end else if (_T_2) begin
        if (_T_3) begin
          if (_T_4) begin
            mem_index <= _T_6;
          end else begin
            mem_index <= _GEN_1;
          end
        end else begin
          mem_index <= _GEN_1;
        end
      end else begin
        mem_index <= _GEN_1;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          mem_data <= odata_hs_io_deq_bits;
        end else if (_T_2) begin
          mem_data <= odata_hs_io_deq_bits;
        end
      end else if (_T_2) begin
        mem_data <= odata_hs_io_deq_bits;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_3) begin
            if (_T_4) begin
              remain <= _T_8;
            end else if (_T_2) begin
              if (_T_3) begin
                if (_T_4) begin
                  remain <= _T_8;
                end else if (_T_1) begin
                  remain <= io_len;
                end
              end else if (_T_1) begin
                remain <= io_len;
              end
            end else if (_T_1) begin
              remain <= io_len;
            end
          end else if (_T_2) begin
            if (_T_3) begin
              if (_T_4) begin
                remain <= _T_8;
              end else if (_T_1) begin
                remain <= io_len;
              end
            end else begin
              remain <= _GEN_3;
            end
          end else begin
            remain <= _GEN_3;
          end
        end else if (_T_2) begin
          if (_T_3) begin
            if (_T_4) begin
              remain <= _T_8;
            end else begin
              remain <= _GEN_3;
            end
          end else begin
            remain <= _GEN_3;
          end
        end else begin
          remain <= _GEN_3;
        end
      end else if (_T_2) begin
        if (_T_3) begin
          if (_T_4) begin
            remain <= _T_8;
          end else begin
            remain <= _GEN_3;
          end
        end else begin
          remain <= _GEN_3;
        end
      end else begin
        remain <= _GEN_3;
      end
    end
  end
endmodule
module LSMemWrapper(
  input         clock,
  input         reset,
  input         io_workEn,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  input         io_readMem_en,
  input  [5:0]  io_readMem_addr,
  output [31:0] io_readMem_dout,
  input         io_writeMem_en,
  input         io_writeMem_we,
  input  [5:0]  io_writeMem_addr,
  input  [31:0] io_writeMem_din,
  input  [5:0]  io_base,
  input  [5:0]  io_len,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits,
  input         io_start,
  input         io_enqEn,
  input         io_deqEn,
  output        io_idle
);
  wire  mem_clock; // @[BasicChiselModules.scala 550:19]
  wire  mem_io_a_en; // @[BasicChiselModules.scala 550:19]
  wire  mem_io_a_we; // @[BasicChiselModules.scala 550:19]
  wire [5:0] mem_io_a_addr; // @[BasicChiselModules.scala 550:19]
  wire [31:0] mem_io_a_din; // @[BasicChiselModules.scala 550:19]
  wire  mem_io_b_en; // @[BasicChiselModules.scala 550:19]
  wire [5:0] mem_io_b_addr; // @[BasicChiselModules.scala 550:19]
  wire [31:0] mem_io_b_dout; // @[BasicChiselModules.scala 550:19]
  wire  enq_mem_clock; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_reset; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_in_ready; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_in_valid; // @[BasicChiselModules.scala 551:23]
  wire [31:0] enq_mem_io_in_bits; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_mem_en; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_mem_we; // @[BasicChiselModules.scala 551:23]
  wire [5:0] enq_mem_io_mem_addr; // @[BasicChiselModules.scala 551:23]
  wire [31:0] enq_mem_io_mem_din; // @[BasicChiselModules.scala 551:23]
  wire [5:0] enq_mem_io_base; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_en; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_start; // @[BasicChiselModules.scala 551:23]
  wire  enq_mem_io_idle; // @[BasicChiselModules.scala 551:23]
  wire  deq_mem_clock; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_reset; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_mem_en; // @[BasicChiselModules.scala 552:23]
  wire [5:0] deq_mem_io_mem_addr; // @[BasicChiselModules.scala 552:23]
  wire [31:0] deq_mem_io_mem_dout; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_out_ready; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_out_valid; // @[BasicChiselModules.scala 552:23]
  wire [31:0] deq_mem_io_out_bits; // @[BasicChiselModules.scala 552:23]
  wire [5:0] deq_mem_io_base; // @[BasicChiselModules.scala 552:23]
  wire [5:0] deq_mem_io_len; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_en; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_start; // @[BasicChiselModules.scala 552:23]
  wire  deq_mem_io_idle; // @[BasicChiselModules.scala 552:23]
  reg [1:0] state; // @[BasicChiselModules.scala 548:22]
  reg [31:0] _RAND_0;
  wire  _T; // @[BasicChiselModules.scala 554:14]
  wire  _GEN_1; // @[BasicChiselModules.scala 559:33]
  wire  _GEN_2; // @[BasicChiselModules.scala 559:33]
  wire [5:0] _GEN_3; // @[BasicChiselModules.scala 559:33]
  wire [31:0] _GEN_4; // @[BasicChiselModules.scala 559:33]
  wire  _GEN_6; // @[BasicChiselModules.scala 555:32]
  wire  _GEN_7; // @[BasicChiselModules.scala 555:32]
  wire [5:0] _GEN_8; // @[BasicChiselModules.scala 555:32]
  wire [31:0] _GEN_9; // @[BasicChiselModules.scala 555:32]
  wire  _T_3; // @[BasicChiselModules.scala 569:20]
  wire  _T_4; // @[BasicChiselModules.scala 570:19]
  wire  _GEN_11; // @[BasicChiselModules.scala 570:32]
  wire  _GEN_12; // @[BasicChiselModules.scala 570:32]
  wire [5:0] _GEN_13; // @[BasicChiselModules.scala 570:32]
  wire [31:0] _GEN_14; // @[BasicChiselModules.scala 570:32]
  wire  _T_5; // @[BasicChiselModules.scala 579:20]
  wire  _GEN_16; // @[BasicChiselModules.scala 580:31]
  wire [5:0] _GEN_17; // @[BasicChiselModules.scala 580:31]
  wire [31:0] _GEN_18; // @[BasicChiselModules.scala 580:31]
  wire  _T_7; // @[BasicChiselModules.scala 591:19]
  wire  _GEN_21; // @[BasicChiselModules.scala 591:32]
  wire [5:0] _GEN_22; // @[BasicChiselModules.scala 591:32]
  wire  _GEN_26; // @[BasicChiselModules.scala 579:32]
  wire [5:0] _GEN_27; // @[BasicChiselModules.scala 579:32]
  wire [31:0] _GEN_28; // @[BasicChiselModules.scala 579:32]
  wire  _GEN_34; // @[BasicChiselModules.scala 579:32]
  wire  _GEN_36; // @[BasicChiselModules.scala 569:38]
  wire  _GEN_37; // @[BasicChiselModules.scala 569:38]
  wire [5:0] _GEN_38; // @[BasicChiselModules.scala 569:38]
  wire [31:0] _GEN_39; // @[BasicChiselModules.scala 569:38]
  wire  _GEN_40; // @[BasicChiselModules.scala 569:38]
  wire [5:0] _GEN_41; // @[BasicChiselModules.scala 569:38]
  wire [31:0] _GEN_42; // @[BasicChiselModules.scala 569:38]
  wire  _GEN_44; // @[BasicChiselModules.scala 569:38]
  SimpleDualPortSram mem ( // @[BasicChiselModules.scala 550:19]
    .clock(mem_clock),
    .io_a_en(mem_io_a_en),
    .io_a_we(mem_io_a_we),
    .io_a_addr(mem_io_a_addr),
    .io_a_din(mem_io_a_din),
    .io_b_en(mem_io_b_en),
    .io_b_addr(mem_io_b_addr),
    .io_b_dout(mem_io_b_dout)
  );
  EnqMem enq_mem ( // @[BasicChiselModules.scala 551:23]
    .clock(enq_mem_clock),
    .reset(enq_mem_reset),
    .io_in_ready(enq_mem_io_in_ready),
    .io_in_valid(enq_mem_io_in_valid),
    .io_in_bits(enq_mem_io_in_bits),
    .io_mem_en(enq_mem_io_mem_en),
    .io_mem_we(enq_mem_io_mem_we),
    .io_mem_addr(enq_mem_io_mem_addr),
    .io_mem_din(enq_mem_io_mem_din),
    .io_base(enq_mem_io_base),
    .io_en(enq_mem_io_en),
    .io_start(enq_mem_io_start),
    .io_idle(enq_mem_io_idle)
  );
  DeqMem deq_mem ( // @[BasicChiselModules.scala 552:23]
    .clock(deq_mem_clock),
    .reset(deq_mem_reset),
    .io_mem_en(deq_mem_io_mem_en),
    .io_mem_addr(deq_mem_io_mem_addr),
    .io_mem_dout(deq_mem_io_mem_dout),
    .io_out_ready(deq_mem_io_out_ready),
    .io_out_valid(deq_mem_io_out_valid),
    .io_out_bits(deq_mem_io_out_bits),
    .io_base(deq_mem_io_base),
    .io_len(deq_mem_io_len),
    .io_en(deq_mem_io_en),
    .io_start(deq_mem_io_start),
    .io_idle(deq_mem_io_idle)
  );
  assign _T = state == 2'h0; // @[BasicChiselModules.scala 554:14]
  assign _GEN_1 = io_enqEn ? enq_mem_io_mem_en : io_writeMem_en; // @[BasicChiselModules.scala 559:33]
  assign _GEN_2 = io_enqEn ? enq_mem_io_mem_we : io_writeMem_we; // @[BasicChiselModules.scala 559:33]
  assign _GEN_3 = io_enqEn ? enq_mem_io_mem_addr : io_writeMem_addr; // @[BasicChiselModules.scala 559:33]
  assign _GEN_4 = io_enqEn ? enq_mem_io_mem_din : io_writeMem_din; // @[BasicChiselModules.scala 559:33]
  assign _GEN_6 = io_workEn ? io_writeMem_en : _GEN_1; // @[BasicChiselModules.scala 555:32]
  assign _GEN_7 = io_workEn ? io_writeMem_we : _GEN_2; // @[BasicChiselModules.scala 555:32]
  assign _GEN_8 = io_workEn ? io_writeMem_addr : _GEN_3; // @[BasicChiselModules.scala 555:32]
  assign _GEN_9 = io_workEn ? io_writeMem_din : _GEN_4; // @[BasicChiselModules.scala 555:32]
  assign _T_3 = state == 2'h1; // @[BasicChiselModules.scala 569:20]
  assign _T_4 = io_enqEn == 1'h0; // @[BasicChiselModules.scala 570:19]
  assign _GEN_11 = _T_4 ? io_writeMem_en : enq_mem_io_mem_en; // @[BasicChiselModules.scala 570:32]
  assign _GEN_12 = _T_4 ? io_writeMem_we : enq_mem_io_mem_we; // @[BasicChiselModules.scala 570:32]
  assign _GEN_13 = _T_4 ? io_writeMem_addr : enq_mem_io_mem_addr; // @[BasicChiselModules.scala 570:32]
  assign _GEN_14 = _T_4 ? io_writeMem_din : enq_mem_io_mem_din; // @[BasicChiselModules.scala 570:32]
  assign _T_5 = state == 2'h2; // @[BasicChiselModules.scala 579:20]
  assign _GEN_16 = io_deqEn ? deq_mem_io_mem_en : io_readMem_en; // @[BasicChiselModules.scala 580:31]
  assign _GEN_17 = io_deqEn ? deq_mem_io_mem_addr : io_readMem_addr; // @[BasicChiselModules.scala 580:31]
  assign _GEN_18 = mem_io_b_dout; // @[BasicChiselModules.scala 580:31]
  assign _T_7 = io_deqEn == 1'h0; // @[BasicChiselModules.scala 591:19]
  assign _GEN_21 = _T_7 ? io_readMem_en : deq_mem_io_mem_en; // @[BasicChiselModules.scala 591:32]
  assign _GEN_22 = _T_7 ? io_readMem_addr : deq_mem_io_mem_addr; // @[BasicChiselModules.scala 591:32]
  assign _GEN_26 = _T_5 ? _GEN_16 : _GEN_21; // @[BasicChiselModules.scala 579:32]
  assign _GEN_27 = _T_5 ? _GEN_17 : _GEN_22; // @[BasicChiselModules.scala 579:32]
  assign _GEN_28 = _T_5 ? _GEN_18 : _GEN_18; // @[BasicChiselModules.scala 579:32]
  assign _GEN_34 = deq_mem_io_idle; // @[BasicChiselModules.scala 579:32]
  assign _GEN_36 = _T_3 ? _GEN_11 : io_writeMem_en; // @[BasicChiselModules.scala 569:38]
  assign _GEN_37 = _T_3 ? _GEN_12 : io_writeMem_we; // @[BasicChiselModules.scala 569:38]
  assign _GEN_38 = _T_3 ? _GEN_13 : io_writeMem_addr; // @[BasicChiselModules.scala 569:38]
  assign _GEN_39 = _T_3 ? _GEN_14 : io_writeMem_din; // @[BasicChiselModules.scala 569:38]
  assign _GEN_40 = _T_3 ? io_readMem_en : _GEN_26; // @[BasicChiselModules.scala 569:38]
  assign _GEN_41 = _T_3 ? io_readMem_addr : _GEN_27; // @[BasicChiselModules.scala 569:38]
  assign _GEN_42 = _T_3 ? mem_io_b_dout : _GEN_28; // @[BasicChiselModules.scala 569:38]
  assign _GEN_44 = _T_3 ? enq_mem_io_idle : _GEN_34; // @[BasicChiselModules.scala 569:38]
  assign io_in_ready = enq_mem_io_in_ready; // @[BasicChiselModules.scala 612:17]
  assign io_readMem_dout = _T ? mem_io_b_dout : _GEN_42; // @[Mem.scala 55:15 Mem.scala 55:15 Mem.scala 55:15 Mem.scala 55:15]
  assign io_out_valid = deq_mem_io_out_valid; // @[BasicChiselModules.scala 616:18]
  assign io_out_bits = deq_mem_io_out_bits; // @[BasicChiselModules.scala 616:18]
  assign io_idle = _T ? enq_mem_io_idle : _GEN_44; // @[BasicChiselModules.scala 568:21 BasicChiselModules.scala 578:21 BasicChiselModules.scala 589:21 BasicChiselModules.scala 600:21]
  assign mem_clock = clock; // @[BasicChiselModules.scala 603:13]
  assign mem_io_a_en = _T ? _GEN_6 : _GEN_36; // @[Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13]
  assign mem_io_a_we = _T ? _GEN_7 : _GEN_37; // @[Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13]
  assign mem_io_a_addr = _T ? _GEN_8 : _GEN_38; // @[Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15]
  assign mem_io_a_din = _T ? _GEN_9 : _GEN_39; // @[Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14]
  assign mem_io_b_en = _T ? io_readMem_en : _GEN_40; // @[Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13]
  assign mem_io_b_addr = _T ? io_readMem_addr : _GEN_41; // @[Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15]
  assign enq_mem_clock = clock; // @[BasicChiselModules.scala 604:17]
  assign enq_mem_reset = reset;
  assign enq_mem_io_in_valid = io_in_valid; // @[BasicChiselModules.scala 612:17]
  assign enq_mem_io_in_bits = io_in_bits; // @[BasicChiselModules.scala 612:17]
  assign enq_mem_io_base = io_base; // @[BasicChiselModules.scala 608:19]
  assign enq_mem_io_en = io_enqEn; // @[BasicChiselModules.scala 611:17]
  assign enq_mem_io_start = io_start; // @[BasicChiselModules.scala 609:20]
  assign deq_mem_clock = clock;
  assign deq_mem_reset = reset;
  assign deq_mem_io_mem_dout = _T_5 ? _GEN_18 : _GEN_18; // @[Mem.scala 55:15 Mem.scala 55:15]
  assign deq_mem_io_out_ready = io_out_ready; // @[BasicChiselModules.scala 616:18]
  assign deq_mem_io_base = io_base; // @[BasicChiselModules.scala 606:19]
  assign deq_mem_io_len = io_len; // @[BasicChiselModules.scala 615:18]
  assign deq_mem_io_en = io_deqEn; // @[BasicChiselModules.scala 614:17]
  assign deq_mem_io_start = io_start; // @[BasicChiselModules.scala 607:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T) begin
      if (io_workEn) begin
        state <= 2'h2;
      end else if (io_enqEn) begin
        state <= 2'h1;
      end
    end else if (_T_3) begin
      if (_T_4) begin
        state <= 2'h2;
      end
    end else if (_T_5) begin
      if (io_deqEn) begin
        state <= 2'h3;
      end
    end else if (_T_7) begin
      state <= 2'h0;
    end
  end
endmodule
module LoadStoreUnit(
  input         clock,
  input         reset,
  input         io_configuration,
  input         io_en,
  input  [3:0]  io_skewing,
  output        io_streamIn_ready,
  input         io_streamIn_valid,
  input  [31:0] io_streamIn_bits,
  input  [5:0]  io_len,
  input         io_streamOut_ready,
  output        io_streamOut_valid,
  output [31:0] io_streamOut_bits,
  input  [5:0]  io_base,
  input         io_start,
  input         io_enqEn,
  input         io_deqEn,
  output        io_idle,
  input  [31:0] io_inputs_1,
  input  [5:0]  io_inputs_0,
  output [31:0] io_outs_0
);
  wire  memWrapper_clock; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_reset; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_workEn; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_in_ready; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_in_valid; // @[BasicChiselModules.scala 645:26]
  wire [31:0] memWrapper_io_in_bits; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_readMem_en; // @[BasicChiselModules.scala 645:26]
  wire [5:0] memWrapper_io_readMem_addr; // @[BasicChiselModules.scala 645:26]
  wire [31:0] memWrapper_io_readMem_dout; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_writeMem_en; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_writeMem_we; // @[BasicChiselModules.scala 645:26]
  wire [5:0] memWrapper_io_writeMem_addr; // @[BasicChiselModules.scala 645:26]
  wire [31:0] memWrapper_io_writeMem_din; // @[BasicChiselModules.scala 645:26]
  wire [5:0] memWrapper_io_base; // @[BasicChiselModules.scala 645:26]
  wire [5:0] memWrapper_io_len; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_out_ready; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_out_valid; // @[BasicChiselModules.scala 645:26]
  wire [31:0] memWrapper_io_out_bits; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_start; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_enqEn; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_deqEn; // @[BasicChiselModules.scala 645:26]
  wire  memWrapper_io_idle; // @[BasicChiselModules.scala 645:26]
  wire  Synchronizer_clock; // @[BasicChiselModules.scala 665:32]
  wire  Synchronizer_reset; // @[BasicChiselModules.scala 665:32]
  wire [3:0] Synchronizer_io_skewing; // @[BasicChiselModules.scala 665:32]
  wire [31:0] Synchronizer_io_input0; // @[BasicChiselModules.scala 665:32]
  wire [31:0] Synchronizer_io_input1; // @[BasicChiselModules.scala 665:32]
  wire [31:0] Synchronizer_io_skewedInput0; // @[BasicChiselModules.scala 665:32]
  wire [31:0] Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 665:32]
  wire  _T; // @[BasicChiselModules.scala 696:27]
  wire  _GEN_1; // @[BasicChiselModules.scala 696:36]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 692:15]
  LSMemWrapper memWrapper ( // @[BasicChiselModules.scala 645:26]
    .clock(memWrapper_clock),
    .reset(memWrapper_reset),
    .io_workEn(memWrapper_io_workEn),
    .io_in_ready(memWrapper_io_in_ready),
    .io_in_valid(memWrapper_io_in_valid),
    .io_in_bits(memWrapper_io_in_bits),
    .io_readMem_en(memWrapper_io_readMem_en),
    .io_readMem_addr(memWrapper_io_readMem_addr),
    .io_readMem_dout(memWrapper_io_readMem_dout),
    .io_writeMem_en(memWrapper_io_writeMem_en),
    .io_writeMem_we(memWrapper_io_writeMem_we),
    .io_writeMem_addr(memWrapper_io_writeMem_addr),
    .io_writeMem_din(memWrapper_io_writeMem_din),
    .io_base(memWrapper_io_base),
    .io_len(memWrapper_io_len),
    .io_out_ready(memWrapper_io_out_ready),
    .io_out_valid(memWrapper_io_out_valid),
    .io_out_bits(memWrapper_io_out_bits),
    .io_start(memWrapper_io_start),
    .io_enqEn(memWrapper_io_enqEn),
    .io_deqEn(memWrapper_io_deqEn),
    .io_idle(memWrapper_io_idle)
  );
  Synchronizer Synchronizer ( // @[BasicChiselModules.scala 665:32]
    .clock(Synchronizer_clock),
    .reset(Synchronizer_reset),
    .io_skewing(Synchronizer_io_skewing),
    .io_input0(Synchronizer_io_input0),
    .io_input1(Synchronizer_io_input1),
    .io_skewedInput0(Synchronizer_io_skewedInput0),
    .io_skewedInput1(Synchronizer_io_skewedInput1)
  );
  assign _T = io_configuration == 1'h0; // @[BasicChiselModules.scala 696:27]
  assign _GEN_1 = _T ? 1'h0 : 1'h1; // @[BasicChiselModules.scala 696:36]
  assign _GEN_2 = Synchronizer_io_skewedInput0; // @[BasicChiselModules.scala 692:15]
  assign io_streamIn_ready = memWrapper_io_in_ready; // @[BasicChiselModules.scala 652:20]
  assign io_streamOut_valid = memWrapper_io_out_valid; // @[BasicChiselModules.scala 653:21]
  assign io_streamOut_bits = memWrapper_io_out_bits; // @[BasicChiselModules.scala 653:21]
  assign io_idle = memWrapper_io_idle; // @[BasicChiselModules.scala 648:22]
  assign io_outs_0 = memWrapper_io_readMem_dout; // @[BasicChiselModules.scala 690:14]
  assign memWrapper_clock = clock;
  assign memWrapper_reset = reset;
  assign memWrapper_io_workEn = io_en; // @[BasicChiselModules.scala 654:24]
  assign memWrapper_io_in_valid = io_streamIn_valid; // @[BasicChiselModules.scala 652:20]
  assign memWrapper_io_in_bits = io_streamIn_bits; // @[BasicChiselModules.scala 652:20]
  assign memWrapper_io_readMem_en = io_en & _T; // @[BasicChiselModules.scala 697:18 BasicChiselModules.scala 701:18 BasicChiselModules.scala 706:16]
  assign memWrapper_io_readMem_addr = _GEN_2[5:0]; // @[BasicChiselModules.scala 693:18]
  assign memWrapper_io_writeMem_en = io_en & _GEN_1; // @[BasicChiselModules.scala 698:19 BasicChiselModules.scala 702:19 BasicChiselModules.scala 707:17]
  assign memWrapper_io_writeMem_we = io_en & _GEN_1; // @[BasicChiselModules.scala 699:19 BasicChiselModules.scala 703:19 BasicChiselModules.scala 708:17]
  assign memWrapper_io_writeMem_addr = _GEN_2[5:0]; // @[BasicChiselModules.scala 694:19]
  assign memWrapper_io_writeMem_din = Synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 695:18]
  assign memWrapper_io_base = io_base; // @[BasicChiselModules.scala 646:22]
  assign memWrapper_io_len = io_len; // @[BasicChiselModules.scala 651:21]
  assign memWrapper_io_out_ready = io_streamOut_ready; // @[BasicChiselModules.scala 653:21]
  assign memWrapper_io_start = io_start; // @[BasicChiselModules.scala 647:23]
  assign memWrapper_io_enqEn = io_enqEn; // @[BasicChiselModules.scala 649:23]
  assign memWrapper_io_deqEn = io_deqEn; // @[BasicChiselModules.scala 650:23]
  assign Synchronizer_clock = clock;
  assign Synchronizer_reset = reset;
  assign Synchronizer_io_skewing = io_skewing; // @[BasicChiselModules.scala 669:31]
  assign Synchronizer_io_input0 = {{26'd0}, io_inputs_0}; // @[BasicChiselModules.scala 666:30]
  assign Synchronizer_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 667:30]
endmodule
module ConfigController(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_II,
  input  [35:0] io_inConfig,
  output [35:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 97:25]
  reg [31:0] _RAND_1;
  reg [35:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_2;
  reg [35:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_3;
  reg [35:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_4;
  reg [35:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_5;
  reg [35:0] configRegs_4; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_6;
  reg [35:0] configRegs_5; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_7;
  reg [35:0] configRegs_6; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_8;
  reg [35:0] configRegs_7; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_9;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [35:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_4; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_5; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_6; // @[BasicChiselModules.scala 106:18]
  wire [35:0] _GEN_7; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [2:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_17; // @[BasicChiselModules.scala 112:32]
  wire [2:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_28; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_38; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 3'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 3'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 3'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _GEN_4 = 3'h4 == cycleReg ? configRegs_4 : _GEN_3; // @[BasicChiselModules.scala 106:18]
  assign _GEN_5 = 3'h5 == cycleReg ? configRegs_5 : _GEN_4; // @[BasicChiselModules.scala 106:18]
  assign _GEN_6 = 3'h6 == cycleReg ? configRegs_6 : _GEN_5; // @[BasicChiselModules.scala 106:18]
  assign _GEN_7 = 3'h7 == cycleReg ? configRegs_7 : _GEN_6; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 3'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_17 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 3'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_28 = _T_1 ? _GEN_17 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_38 = io_en & _GEN_28; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 36'h0 : _GEN_7; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  configRegs_0 = _RAND_2[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  configRegs_1 = _RAND_3[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  configRegs_2 = _RAND_4[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  configRegs_3 = _RAND_5[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  configRegs_4 = _RAND_6[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  configRegs_5 = _RAND_7[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  configRegs_6 = _RAND_8[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  configRegs_7 = _RAND_9[35:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_38;
    end
    if (reset) begin
      cycleReg <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 3'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 3'h0;
    end
    if (reset) begin
      configRegs_0 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_4 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h4 == cycleReg) begin
          configRegs_4 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_5 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h5 == cycleReg) begin
          configRegs_5 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_6 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h6 == cycleReg) begin
          configRegs_6 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_7 <= 36'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h7 == cycleReg) begin
          configRegs_7 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_145(
  input  [35:0] io_configuration,
  output [2:0]  io_outs_11,
  output [2:0]  io_outs_10,
  output [2:0]  io_outs_9,
  output [2:0]  io_outs_8,
  output [2:0]  io_outs_7,
  output [2:0]  io_outs_6,
  output [2:0]  io_outs_5,
  output [2:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [2:0]  io_outs_0
);
  assign io_outs_11 = io_configuration[35:33]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_10 = io_configuration[32:30]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_9 = io_configuration[29:27]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_8 = io_configuration[26:24]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_7 = io_configuration[23:21]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_6 = io_configuration[20:18]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_5 = io_configuration[17:15]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_4 = io_configuration[14:12]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_3 = io_configuration[11:9]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_2 = io_configuration[8:6]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_1 = io_configuration[5:3]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[2:0]; // @[BasicChiselModules.scala 490:18]
endmodule
module ConfigController_2(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_II,
  input  [59:0] io_inConfig,
  output [59:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 97:25]
  reg [31:0] _RAND_1;
  reg [59:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_2;
  reg [59:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_3;
  reg [59:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_4;
  reg [59:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_5;
  reg [59:0] configRegs_4; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_6;
  reg [59:0] configRegs_5; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_7;
  reg [59:0] configRegs_6; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_8;
  reg [59:0] configRegs_7; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_9;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [59:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_4; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_5; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_6; // @[BasicChiselModules.scala 106:18]
  wire [59:0] _GEN_7; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [2:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_17; // @[BasicChiselModules.scala 112:32]
  wire [2:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_28; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_38; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 3'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 3'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 3'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _GEN_4 = 3'h4 == cycleReg ? configRegs_4 : _GEN_3; // @[BasicChiselModules.scala 106:18]
  assign _GEN_5 = 3'h5 == cycleReg ? configRegs_5 : _GEN_4; // @[BasicChiselModules.scala 106:18]
  assign _GEN_6 = 3'h6 == cycleReg ? configRegs_6 : _GEN_5; // @[BasicChiselModules.scala 106:18]
  assign _GEN_7 = 3'h7 == cycleReg ? configRegs_7 : _GEN_6; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 3'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_17 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 3'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_28 = _T_1 ? _GEN_17 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_38 = io_en & _GEN_28; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 60'h0 : _GEN_7; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  configRegs_0 = _RAND_2[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  configRegs_1 = _RAND_3[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  configRegs_2 = _RAND_4[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  configRegs_3 = _RAND_5[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  configRegs_4 = _RAND_6[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  configRegs_5 = _RAND_7[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  configRegs_6 = _RAND_8[59:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  configRegs_7 = _RAND_9[59:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_38;
    end
    if (reset) begin
      cycleReg <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 3'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 3'h0;
    end
    if (reset) begin
      configRegs_0 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_4 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h4 == cycleReg) begin
          configRegs_4 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_5 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h5 == cycleReg) begin
          configRegs_5 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_6 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h6 == cycleReg) begin
          configRegs_6 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_7 <= 60'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h7 == cycleReg) begin
          configRegs_7 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_147(
  input  [59:0] io_configuration,
  output        io_outs_12,
  output [31:0] io_outs_11,
  output        io_outs_10,
  output        io_outs_9,
  output        io_outs_8,
  output [2:0]  io_outs_7,
  output [2:0]  io_outs_6,
  output [2:0]  io_outs_5,
  output [2:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [2:0]  io_outs_0
);
  assign io_outs_12 = io_configuration[59]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_11 = io_configuration[58:27]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_10 = io_configuration[26]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_9 = io_configuration[25]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_8 = io_configuration[24]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_7 = io_configuration[23:21]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_6 = io_configuration[20:18]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_5 = io_configuration[17:15]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_4 = io_configuration[14:12]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_3 = io_configuration[11:9]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_2 = io_configuration[8:6]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_1 = io_configuration[5:3]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[2:0]; // @[BasicChiselModules.scala 490:18]
endmodule
module ConfigController_3(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_II,
  input  [75:0] io_inConfig,
  output [75:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 97:25]
  reg [31:0] _RAND_1;
  reg [75:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_2;
  reg [75:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_3;
  reg [75:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_4;
  reg [75:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_5;
  reg [75:0] configRegs_4; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_6;
  reg [75:0] configRegs_5; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_7;
  reg [75:0] configRegs_6; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_8;
  reg [75:0] configRegs_7; // @[BasicChiselModules.scala 99:27]
  reg [95:0] _RAND_9;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [75:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_4; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_5; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_6; // @[BasicChiselModules.scala 106:18]
  wire [75:0] _GEN_7; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [2:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_17; // @[BasicChiselModules.scala 112:32]
  wire [2:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_28; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_38; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 3'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 3'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 3'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _GEN_4 = 3'h4 == cycleReg ? configRegs_4 : _GEN_3; // @[BasicChiselModules.scala 106:18]
  assign _GEN_5 = 3'h5 == cycleReg ? configRegs_5 : _GEN_4; // @[BasicChiselModules.scala 106:18]
  assign _GEN_6 = 3'h6 == cycleReg ? configRegs_6 : _GEN_5; // @[BasicChiselModules.scala 106:18]
  assign _GEN_7 = 3'h7 == cycleReg ? configRegs_7 : _GEN_6; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 3'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_17 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 3'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_28 = _T_1 ? _GEN_17 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_38 = io_en & _GEN_28; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 76'h0 : _GEN_7; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {3{`RANDOM}};
  configRegs_0 = _RAND_2[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  configRegs_1 = _RAND_3[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {3{`RANDOM}};
  configRegs_2 = _RAND_4[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  configRegs_3 = _RAND_5[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  configRegs_4 = _RAND_6[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  configRegs_5 = _RAND_7[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {3{`RANDOM}};
  configRegs_6 = _RAND_8[75:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {3{`RANDOM}};
  configRegs_7 = _RAND_9[75:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_38;
    end
    if (reset) begin
      cycleReg <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 3'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 3'h0;
    end
    if (reset) begin
      configRegs_0 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_4 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h4 == cycleReg) begin
          configRegs_4 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_5 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h5 == cycleReg) begin
          configRegs_5 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_6 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h6 == cycleReg) begin
          configRegs_6 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_7 <= 76'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h7 == cycleReg) begin
          configRegs_7 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_148(
  input  [75:0] io_configuration,
  output [31:0] io_outs_17,
  output        io_outs_16,
  output        io_outs_15,
  output        io_outs_14,
  output        io_outs_13,
  output [2:0]  io_outs_12,
  output [2:0]  io_outs_11,
  output [2:0]  io_outs_10,
  output [2:0]  io_outs_9,
  output [2:0]  io_outs_8,
  output [2:0]  io_outs_7,
  output [2:0]  io_outs_6,
  output [2:0]  io_outs_5,
  output [2:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [3:0]  io_outs_0
);
  assign io_outs_17 = io_configuration[75:44]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_16 = io_configuration[43]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_15 = io_configuration[42]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_14 = io_configuration[41]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_13 = io_configuration[40]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_12 = io_configuration[39:37]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_11 = io_configuration[36:34]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_10 = io_configuration[33:31]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_9 = io_configuration[30:28]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_8 = io_configuration[27:25]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_7 = io_configuration[24:22]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_6 = io_configuration[21:19]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_5 = io_configuration[18:16]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_4 = io_configuration[15:13]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_3 = io_configuration[12:10]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_2 = io_configuration[9:7]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_1 = io_configuration[6:4]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[3:0]; // @[BasicChiselModules.scala 490:18]
endmodule
module Dispatch_171(
  input  [1767:0] io_configuration,
  output [59:0]   io_outs_25,
  output [75:0]   io_outs_24,
  output [75:0]   io_outs_23,
  output [75:0]   io_outs_22,
  output [75:0]   io_outs_21,
  output [59:0]   io_outs_20,
  output [59:0]   io_outs_19,
  output [75:0]   io_outs_18,
  output [75:0]   io_outs_17,
  output [75:0]   io_outs_16,
  output [75:0]   io_outs_15,
  output [59:0]   io_outs_14,
  output [59:0]   io_outs_13,
  output [75:0]   io_outs_12,
  output [75:0]   io_outs_11,
  output [75:0]   io_outs_10,
  output [75:0]   io_outs_9,
  output [59:0]   io_outs_8,
  output [59:0]   io_outs_7,
  output [75:0]   io_outs_6,
  output [75:0]   io_outs_5,
  output [75:0]   io_outs_4,
  output [75:0]   io_outs_3,
  output [59:0]   io_outs_2,
  output [35:0]   io_outs_1,
  output [35:0]   io_outs_0
);
  assign io_outs_25 = io_configuration[1767:1708]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_24 = io_configuration[1707:1632]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_23 = io_configuration[1631:1556]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_22 = io_configuration[1555:1480]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_21 = io_configuration[1479:1404]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_20 = io_configuration[1403:1344]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_19 = io_configuration[1343:1284]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_18 = io_configuration[1283:1208]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_17 = io_configuration[1207:1132]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_16 = io_configuration[1131:1056]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_15 = io_configuration[1055:980]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_14 = io_configuration[979:920]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_13 = io_configuration[919:860]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_12 = io_configuration[859:784]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_11 = io_configuration[783:708]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_10 = io_configuration[707:632]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_9 = io_configuration[631:556]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_8 = io_configuration[555:496]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_7 = io_configuration[495:436]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_6 = io_configuration[435:360]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_5 = io_configuration[359:284]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_4 = io_configuration[283:208]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_3 = io_configuration[207:132]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_2 = io_configuration[131:72]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_1 = io_configuration[71:36]; // @[BasicChiselModules.scala 490:18]
  assign io_outs_0 = io_configuration[35:0]; // @[BasicChiselModules.scala 490:18]
endmodule
module TopModule(
  input           clock,
  input           reset,
  output          io_streamInLSU_7_ready,
  input           io_streamInLSU_7_valid,
  input  [31:0]   io_streamInLSU_7_bits,
  output          io_streamInLSU_6_ready,
  input           io_streamInLSU_6_valid,
  input  [31:0]   io_streamInLSU_6_bits,
  output          io_streamInLSU_5_ready,
  input           io_streamInLSU_5_valid,
  input  [31:0]   io_streamInLSU_5_bits,
  output          io_streamInLSU_4_ready,
  input           io_streamInLSU_4_valid,
  input  [31:0]   io_streamInLSU_4_bits,
  output          io_streamInLSU_3_ready,
  input           io_streamInLSU_3_valid,
  input  [31:0]   io_streamInLSU_3_bits,
  output          io_streamInLSU_2_ready,
  input           io_streamInLSU_2_valid,
  input  [31:0]   io_streamInLSU_2_bits,
  output          io_streamInLSU_1_ready,
  input           io_streamInLSU_1_valid,
  input  [31:0]   io_streamInLSU_1_bits,
  output          io_streamInLSU_0_ready,
  input           io_streamInLSU_0_valid,
  input  [31:0]   io_streamInLSU_0_bits,
  input           io_streamOutLSU_7_ready,
  output          io_streamOutLSU_7_valid,
  output [31:0]   io_streamOutLSU_7_bits,
  input           io_streamOutLSU_6_ready,
  output          io_streamOutLSU_6_valid,
  output [31:0]   io_streamOutLSU_6_bits,
  input           io_streamOutLSU_5_ready,
  output          io_streamOutLSU_5_valid,
  output [31:0]   io_streamOutLSU_5_bits,
  input           io_streamOutLSU_4_ready,
  output          io_streamOutLSU_4_valid,
  output [31:0]   io_streamOutLSU_4_bits,
  input           io_streamOutLSU_3_ready,
  output          io_streamOutLSU_3_valid,
  output [31:0]   io_streamOutLSU_3_bits,
  input           io_streamOutLSU_2_ready,
  output          io_streamOutLSU_2_valid,
  output [31:0]   io_streamOutLSU_2_bits,
  input           io_streamOutLSU_1_ready,
  output          io_streamOutLSU_1_valid,
  output [31:0]   io_streamOutLSU_1_bits,
  input           io_streamOutLSU_0_ready,
  output          io_streamOutLSU_0_valid,
  output [31:0]   io_streamOutLSU_0_bits,
  input  [5:0]    io_baseLSU_0,
  input  [5:0]    io_baseLSU_1,
  input  [5:0]    io_baseLSU_2,
  input  [5:0]    io_baseLSU_3,
  input  [5:0]    io_baseLSU_4,
  input  [5:0]    io_baseLSU_5,
  input  [5:0]    io_baseLSU_6,
  input  [5:0]    io_baseLSU_7,
  input  [5:0]    io_lenLSU_0,
  input  [5:0]    io_lenLSU_1,
  input  [5:0]    io_lenLSU_2,
  input  [5:0]    io_lenLSU_3,
  input  [5:0]    io_lenLSU_4,
  input  [5:0]    io_lenLSU_5,
  input  [5:0]    io_lenLSU_6,
  input  [5:0]    io_lenLSU_7,
  input           io_startLSU_0,
  input           io_startLSU_1,
  input           io_startLSU_2,
  input           io_startLSU_3,
  input           io_startLSU_4,
  input           io_startLSU_5,
  input           io_startLSU_6,
  input           io_startLSU_7,
  input           io_enqEnLSU_0,
  input           io_enqEnLSU_1,
  input           io_enqEnLSU_2,
  input           io_enqEnLSU_3,
  input           io_enqEnLSU_4,
  input           io_enqEnLSU_5,
  input           io_enqEnLSU_6,
  input           io_enqEnLSU_7,
  input           io_deqEnLSU_0,
  input           io_deqEnLSU_1,
  input           io_deqEnLSU_2,
  input           io_deqEnLSU_3,
  input           io_deqEnLSU_4,
  input           io_deqEnLSU_5,
  input           io_deqEnLSU_6,
  input           io_deqEnLSU_7,
  output          io_idleLSU_0,
  output          io_idleLSU_1,
  output          io_idleLSU_2,
  output          io_idleLSU_3,
  output          io_idleLSU_4,
  output          io_idleLSU_5,
  output          io_idleLSU_6,
  output          io_idleLSU_7,
  input           io_enConfig,
  input           io_en,
  input  [1151:0] io_schedules,
  input  [2:0]    io_II,
  input  [1767:0] io_configuration,
  input  [31:0]   io_inputs_11,
  input  [31:0]   io_inputs_10,
  input  [31:0]   io_inputs_9,
  input  [31:0]   io_inputs_8,
  input  [31:0]   io_inputs_7,
  input  [31:0]   io_inputs_6,
  input  [31:0]   io_inputs_5,
  input  [31:0]   io_inputs_4,
  input  [31:0]   io_inputs_3,
  input  [31:0]   io_inputs_2,
  input  [31:0]   io_inputs_1,
  input  [31:0]   io_inputs_0,
  output [31:0]   io_outs_11,
  output [31:0]   io_outs_10,
  output [31:0]   io_outs_9,
  output [31:0]   io_outs_8,
  output [31:0]   io_outs_7,
  output [31:0]   io_outs_6,
  output [31:0]   io_outs_5,
  output [31:0]   io_outs_4,
  output [31:0]   io_outs_3,
  output [31:0]   io_outs_2,
  output [31:0]   io_outs_1,
  output [31:0]   io_outs_0
);
  wire [1151:0] Dispatch_io_configuration; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_191; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_190; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_189; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_188; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_187; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_186; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_185; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_184; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_183; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_182; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_181; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_180; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_179; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_178; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_177; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_176; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_175; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_174; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_173; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_172; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_171; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_170; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_169; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_168; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_167; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_166; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_165; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_164; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_163; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_162; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_161; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_160; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_159; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_158; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_157; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_156; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_155; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_154; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_153; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_152; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_151; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_150; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_149; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_148; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_147; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_146; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_145; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_144; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_143; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_142; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_141; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_140; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_139; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_138; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_137; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_136; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_135; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_134; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_133; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_132; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_131; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_130; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_129; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_128; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_127; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_126; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_125; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_124; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_123; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_122; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_121; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_120; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_119; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_118; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_117; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_116; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_115; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_114; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_113; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_112; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_111; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_110; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_109; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_108; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_107; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_106; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_105; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_104; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_103; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_102; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_101; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_100; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_99; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_98; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_97; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_96; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_95; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_94; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_93; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_92; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_91; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_90; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_89; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_88; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_87; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_86; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_85; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_84; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_83; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_82; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_81; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_80; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_79; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_78; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_77; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_76; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_75; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_74; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_73; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_72; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_71; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_70; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_69; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_68; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_67; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_66; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_65; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_64; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_63; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_62; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_61; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_60; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_59; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_58; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_57; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_56; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_55; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_54; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_53; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_52; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_51; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_50; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_49; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_48; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_47; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_46; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_45; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_44; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_43; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_42; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_41; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_40; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_39; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_38; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_37; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_36; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_35; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_34; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_33; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_32; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_31; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_30; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_29; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_28; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_27; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_26; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_25; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_24; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_23; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_22; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_21; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_20; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_19; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_18; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_17; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_16; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_15; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_14; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_13; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_12; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_11; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_10; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_9; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_8; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_7; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_6; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_5; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_4; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_3; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_2; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_1; // @[TopModule.scala 122:34]
  wire [5:0] Dispatch_io_outs_0; // @[TopModule.scala 122:34]
  wire  Alu_clock; // @[TopModule.scala 131:54]
  wire  Alu_reset; // @[TopModule.scala 131:54]
  wire  Alu_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_1_clock; // @[TopModule.scala 131:54]
  wire  Alu_1_reset; // @[TopModule.scala 131:54]
  wire  Alu_1_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_1_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_1_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_1_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_1_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_1_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_2_clock; // @[TopModule.scala 131:54]
  wire  Alu_2_reset; // @[TopModule.scala 131:54]
  wire  Alu_2_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_2_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_2_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_2_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_2_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_2_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_3_clock; // @[TopModule.scala 131:54]
  wire  Alu_3_reset; // @[TopModule.scala 131:54]
  wire  Alu_3_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_3_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_3_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_3_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_3_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_3_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_4_clock; // @[TopModule.scala 131:54]
  wire  Alu_4_reset; // @[TopModule.scala 131:54]
  wire  Alu_4_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_4_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_4_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_4_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_4_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_4_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_5_clock; // @[TopModule.scala 131:54]
  wire  Alu_5_reset; // @[TopModule.scala 131:54]
  wire  Alu_5_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_5_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_5_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_5_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_5_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_5_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_6_clock; // @[TopModule.scala 131:54]
  wire  Alu_6_reset; // @[TopModule.scala 131:54]
  wire  Alu_6_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_6_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_6_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_6_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_6_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_6_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_7_clock; // @[TopModule.scala 131:54]
  wire  Alu_7_reset; // @[TopModule.scala 131:54]
  wire  Alu_7_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_7_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_7_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_7_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_7_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_7_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_8_clock; // @[TopModule.scala 131:54]
  wire  Alu_8_reset; // @[TopModule.scala 131:54]
  wire  Alu_8_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_8_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_8_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_8_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_8_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_8_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_9_clock; // @[TopModule.scala 131:54]
  wire  Alu_9_reset; // @[TopModule.scala 131:54]
  wire  Alu_9_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_9_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_9_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_9_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_9_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_9_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_10_clock; // @[TopModule.scala 131:54]
  wire  Alu_10_reset; // @[TopModule.scala 131:54]
  wire  Alu_10_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_10_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_10_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_10_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_10_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_10_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_11_clock; // @[TopModule.scala 131:54]
  wire  Alu_11_reset; // @[TopModule.scala 131:54]
  wire  Alu_11_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_11_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_11_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_11_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_11_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_11_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_12_clock; // @[TopModule.scala 131:54]
  wire  Alu_12_reset; // @[TopModule.scala 131:54]
  wire  Alu_12_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_12_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_12_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_12_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_12_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_12_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_13_clock; // @[TopModule.scala 131:54]
  wire  Alu_13_reset; // @[TopModule.scala 131:54]
  wire  Alu_13_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_13_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_13_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_13_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_13_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_13_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_14_clock; // @[TopModule.scala 131:54]
  wire  Alu_14_reset; // @[TopModule.scala 131:54]
  wire  Alu_14_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_14_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_14_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_14_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_14_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_14_io_outs_0; // @[TopModule.scala 131:54]
  wire  Alu_15_clock; // @[TopModule.scala 131:54]
  wire  Alu_15_reset; // @[TopModule.scala 131:54]
  wire  Alu_15_io_en; // @[TopModule.scala 131:54]
  wire [3:0] Alu_15_io_skewing; // @[TopModule.scala 131:54]
  wire [3:0] Alu_15_io_configuration; // @[TopModule.scala 131:54]
  wire [31:0] Alu_15_io_inputs_1; // @[TopModule.scala 131:54]
  wire [31:0] Alu_15_io_inputs_0; // @[TopModule.scala 131:54]
  wire [31:0] Alu_15_io_outs_0; // @[TopModule.scala 131:54]
  wire  MultiIIScheduleController_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_1_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_1_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_1_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_1_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_1_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_1_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_2_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_2_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_2_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_2_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_2_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_2_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_3_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_3_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_3_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_3_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_3_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_3_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_4_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_4_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_4_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_4_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_4_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_4_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_5_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_5_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_5_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_5_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_5_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_5_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_6_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_6_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_6_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_6_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_6_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_6_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_7_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_7_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_7_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_7_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_7_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_7_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_8_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_8_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_8_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_8_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_8_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_8_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_9_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_9_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_9_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_9_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_9_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_9_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_10_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_10_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_10_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_10_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_10_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_10_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_11_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_11_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_11_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_11_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_11_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_11_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_12_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_12_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_12_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_12_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_12_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_12_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_13_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_13_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_13_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_13_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_13_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_13_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_14_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_14_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_14_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_14_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_14_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_14_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_15_clock; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_15_reset; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_15_io_en; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_0; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_1; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_2; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_3; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_4; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_5; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_6; // @[TopModule.scala 135:23]
  wire [5:0] MultiIIScheduleController_15_io_schedules_7; // @[TopModule.scala 135:23]
  wire [2:0] MultiIIScheduleController_15_io_II; // @[TopModule.scala 135:23]
  wire  MultiIIScheduleController_15_io_valid; // @[TopModule.scala 135:23]
  wire [3:0] MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 135:23]
  wire  RegisterFile_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_1_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_1_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_1_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_1_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_1_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_2_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_2_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_2_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_2_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_2_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_3_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_3_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_3_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_3_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_3_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_4_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_4_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_4_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_4_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_4_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_5_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_5_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_5_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_5_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_5_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_6_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_6_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_6_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_6_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_6_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_7_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_7_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_7_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_7_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_7_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_8_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_8_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_8_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_8_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_8_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_9_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_9_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_9_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_9_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_9_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_10_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_10_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_10_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_10_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_10_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_11_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_11_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_11_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_11_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_11_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_12_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_12_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_12_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_12_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_12_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_13_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_13_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_13_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_13_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_13_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_14_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_14_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_14_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_14_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_14_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_15_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_15_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_15_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_15_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_15_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_16_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_16_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_16_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_16_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_16_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_17_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_17_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_17_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_17_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_17_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_18_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_18_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_18_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_18_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_18_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_19_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_19_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_19_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_19_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_19_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_20_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_20_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_20_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_20_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_20_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_21_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_21_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_21_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_21_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_21_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_22_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_22_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_22_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_22_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_22_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_23_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_23_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_23_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_23_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_23_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_24_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_24_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_24_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_24_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_24_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_25_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_25_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_25_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_25_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_25_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_26_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_26_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_26_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_26_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_26_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_27_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_27_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_27_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_27_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_27_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_28_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_28_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_28_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_28_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_28_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_29_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_29_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_29_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_29_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_29_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_30_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_30_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_30_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_30_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_30_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_31_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_31_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_31_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_31_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_31_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_32_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_32_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_32_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_32_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_32_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_33_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_33_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_33_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_33_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_33_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_34_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_34_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_34_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_34_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_34_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_35_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_35_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_35_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_35_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_35_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_36_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_36_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_36_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_36_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_36_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_37_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_37_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_37_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_37_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_37_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_38_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_38_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_38_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_38_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_38_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_39_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_39_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_39_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_39_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_39_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_40_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_40_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_40_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_40_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_40_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_41_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_41_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_41_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_41_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_41_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_42_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_42_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_42_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_42_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_42_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_43_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_43_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_43_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_43_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_43_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_44_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_44_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_44_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_44_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_44_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_45_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_45_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_45_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_45_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_45_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_46_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_46_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_46_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_46_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_46_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_47_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_47_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_47_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_47_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_47_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_48_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_48_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_48_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_48_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_48_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_49_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_49_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_49_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_49_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_49_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_50_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_50_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_50_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_50_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_50_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_51_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_51_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_51_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_51_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_51_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_52_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_52_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_52_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_52_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_52_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_53_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_53_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_53_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_53_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_53_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_54_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_54_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_54_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_54_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_54_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_55_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_55_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_55_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_55_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_55_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_56_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_56_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_56_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_56_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_56_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_57_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_57_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_57_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_57_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_57_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_58_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_58_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_58_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_58_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_58_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_59_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_59_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_59_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_59_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_59_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_60_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_60_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_60_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_60_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_60_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_61_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_61_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_61_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_61_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_61_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_62_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_62_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_62_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_62_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_62_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_63_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_63_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_63_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_63_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_63_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_64_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_64_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_64_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_64_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_64_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_65_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_65_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_65_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_65_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_65_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_66_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_66_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_66_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_66_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_66_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_67_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_67_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_67_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_67_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_67_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_68_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_68_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_68_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_68_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_68_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_69_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_69_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_69_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_69_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_69_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_70_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_70_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_70_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_70_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_70_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_71_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_71_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_71_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_71_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_71_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_72_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_72_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_72_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_72_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_72_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_73_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_73_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_73_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_73_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_73_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_74_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_74_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_74_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_74_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_74_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_75_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_75_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_75_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_75_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_75_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_76_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_76_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_76_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_76_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_76_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_77_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_77_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_77_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_77_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_77_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_78_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_78_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_78_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_78_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_78_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_79_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_79_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_79_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_79_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_79_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_80_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_80_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_80_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_80_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_80_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_81_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_81_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_81_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_81_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_81_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_82_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_82_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_82_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_82_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_82_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_83_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_83_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_83_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_83_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_83_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_84_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_84_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_84_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_84_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_84_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_85_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_85_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_85_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_85_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_85_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_86_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_86_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_86_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_86_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_86_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_87_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_87_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_87_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_87_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_87_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_88_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_88_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_88_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_88_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_88_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_89_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_89_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_89_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_89_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_89_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_90_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_90_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_90_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_90_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_90_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_91_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_91_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_91_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_91_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_91_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_92_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_92_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_92_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_92_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_92_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_93_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_93_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_93_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_93_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_93_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_94_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_94_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_94_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_94_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_94_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_95_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_95_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_95_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_95_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_95_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_96_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_96_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_96_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_96_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_96_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_97_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_97_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_97_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_97_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_97_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_98_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_98_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_98_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_98_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_98_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_99_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_99_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_99_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_99_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_99_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_100_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_100_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_100_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_100_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_100_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_101_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_101_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_101_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_101_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_101_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_102_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_102_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_102_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_102_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_102_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_103_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_103_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_103_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_103_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_103_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_104_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_104_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_104_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_104_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_104_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_105_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_105_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_105_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_105_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_105_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_106_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_106_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_106_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_106_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_106_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_107_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_107_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_107_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_107_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_107_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_108_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_108_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_108_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_108_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_108_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_109_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_109_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_109_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_109_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_109_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_110_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_110_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_110_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_110_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_110_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_111_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_111_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_111_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_111_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_111_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_112_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_112_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_112_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_112_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_112_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_113_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_113_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_113_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_113_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_113_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_114_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_114_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_114_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_114_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_114_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_115_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_115_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_115_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_115_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_115_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_116_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_116_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_116_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_116_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_116_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_117_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_117_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_117_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_117_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_117_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_118_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_118_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_118_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_118_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_118_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_119_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_119_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_119_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_119_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_119_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_120_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_120_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_120_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_120_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_120_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_121_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_121_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_121_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_121_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_121_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_122_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_122_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_122_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_122_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_122_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_123_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_123_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_123_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_123_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_123_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_124_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_124_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_124_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_124_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_124_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_125_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_125_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_125_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_125_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_125_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_126_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_126_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_126_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_126_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_126_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_127_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_127_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_127_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_127_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_127_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_128_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_128_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_128_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_128_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_128_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_129_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_129_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_129_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_129_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_129_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_130_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_130_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_130_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_130_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_130_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_131_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_131_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_131_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_131_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_131_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_132_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_132_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_132_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_132_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_132_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_133_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_133_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_133_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_133_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_133_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_134_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_134_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_134_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_134_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_134_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_135_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_135_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_135_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_135_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_135_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_136_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_136_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_136_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_136_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_136_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_137_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_137_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_137_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_137_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_137_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_138_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_138_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_138_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_138_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_138_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_139_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_139_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_139_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_139_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_139_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_140_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_140_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_140_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_140_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_140_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_141_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_141_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_141_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_141_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_141_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_142_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_142_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_142_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_142_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_142_io_outs_0; // @[TopModule.scala 158:21]
  wire  RegisterFile_143_clock; // @[TopModule.scala 158:21]
  wire  RegisterFile_143_reset; // @[TopModule.scala 158:21]
  wire [2:0] RegisterFile_143_io_configuration; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_143_io_inputs_0; // @[TopModule.scala 158:21]
  wire [31:0] RegisterFile_143_io_outs_0; // @[TopModule.scala 158:21]
  wire [2:0] Multiplexer_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_1_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_1_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_2_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_2_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_3_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_3_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_4_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_4_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_5_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_5_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_5_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_5_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_6_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_6_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_6_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_6_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_7_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_7_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_7_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_7_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_8_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_8_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_9_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_9_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_10_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_10_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_11_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_11_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_12_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_12_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_13_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_13_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_14_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_14_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_14_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_14_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_15_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_15_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_15_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_15_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_16_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_16_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_16_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_16_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_17_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_17_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_17_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_17_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_18_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_18_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_19_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_19_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_20_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_20_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_21_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_21_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_22_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_22_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_23_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_23_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_24_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_24_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_24_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_24_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_25_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_25_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_25_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_25_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_26_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_26_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_26_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_26_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_27_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_27_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_27_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_27_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_28_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_28_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_29_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_29_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_30_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_30_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_31_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_31_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_32_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_32_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_33_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_33_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_34_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_34_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_34_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_34_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_35_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_35_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_35_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_35_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_36_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_36_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_36_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_36_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_37_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_37_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_37_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_37_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_38_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_38_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_39_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_39_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_40_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_40_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_41_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_41_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_42_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_42_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_43_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_43_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_44_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_44_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_44_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_44_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_45_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_45_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_45_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_45_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_46_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_46_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_46_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_46_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_47_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_47_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_47_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_47_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_48_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_48_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_49_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_49_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_50_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_50_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_51_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_51_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_52_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_52_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_53_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_53_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_53_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_53_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_54_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_54_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_54_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_54_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_55_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_55_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_55_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_55_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_56_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_56_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_57_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_57_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_58_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_58_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_59_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_59_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_60_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_60_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_61_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_61_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_61_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_61_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_62_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_62_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_62_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_62_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_63_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_63_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_63_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_63_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_64_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_64_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_65_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_65_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_66_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_66_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_67_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_67_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_68_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_68_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_69_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_69_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_70_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_70_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_70_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_70_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_71_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_71_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_71_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_71_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_72_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_72_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_72_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_72_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_73_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_73_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_73_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_73_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_74_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_74_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_75_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_75_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_76_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_76_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_77_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_77_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_78_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_78_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_79_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_79_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_80_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_80_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_80_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_80_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_81_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_81_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_81_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_81_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_82_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_82_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_82_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_82_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_83_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_83_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_83_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_83_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_84_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_84_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_85_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_85_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_86_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_86_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_87_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_87_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_88_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_88_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_89_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_89_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_90_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_90_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_90_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_90_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_91_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_91_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_91_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_91_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_92_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_92_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_92_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_92_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_93_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_93_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_93_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_93_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_94_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_94_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_95_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_95_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_96_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_96_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_97_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_97_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_98_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_98_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_99_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_99_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_100_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_100_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_100_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_100_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_101_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_101_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_101_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_101_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_102_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_102_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_102_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_102_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_103_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_103_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_103_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_103_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_104_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_104_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_105_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_105_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_106_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_106_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_107_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_107_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_108_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_108_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_109_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_109_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_109_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_109_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_110_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_110_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_110_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_110_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_111_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_111_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_111_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_111_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_112_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_112_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_113_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_113_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_114_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_114_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_115_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_115_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_116_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_116_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_117_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_117_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_117_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_117_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_118_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_118_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_118_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_118_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_119_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_119_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_119_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_119_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_120_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_120_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_121_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_121_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_122_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_122_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_123_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_123_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_124_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_124_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_125_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_125_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_126_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_126_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_126_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_126_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_127_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_127_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_127_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_127_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_128_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_128_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_128_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_128_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_129_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_129_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_129_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_129_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_130_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_130_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_131_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_131_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_132_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_132_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_133_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_133_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_134_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_134_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_135_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_135_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_136_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_136_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_136_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_136_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_137_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_137_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_137_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_137_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_138_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_138_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_138_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_138_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_139_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_139_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_139_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_139_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_140_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_140_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_141_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_141_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_142_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_142_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_143_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_143_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_144_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_144_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_145_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_145_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_146_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_146_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_146_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_146_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_147_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_147_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_147_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_147_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_148_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_148_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_148_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_148_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_149_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_149_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_149_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_149_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_150_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_150_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_151_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_151_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_152_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_152_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_153_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_153_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_154_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_154_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_155_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_155_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_156_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_156_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_156_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_156_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_157_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_157_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_157_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_157_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_158_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_158_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_158_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_158_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_159_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_159_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_159_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_159_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_160_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_160_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_161_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_161_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_162_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_162_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_163_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_163_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_164_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_164_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_165_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_165_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_165_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_165_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_166_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_166_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_166_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_166_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_167_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_167_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_167_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_167_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_168_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_168_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_169_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_169_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_170_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_170_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_171_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_171_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_172_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_172_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_173_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_173_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_173_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_173_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_174_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_174_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_174_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_174_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_175_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_175_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_175_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_175_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_176_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_176_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_177_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_177_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_178_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_178_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_179_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_179_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_180_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_180_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_181_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_181_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_182_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_182_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_182_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_182_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_183_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_183_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_183_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_183_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_184_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_184_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_184_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_184_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_185_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_185_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_185_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_185_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_186_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_186_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_187_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_187_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_188_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_188_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_189_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_189_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_190_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_190_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_191_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_191_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_192_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_192_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_192_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_192_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_193_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_193_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_193_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_193_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_194_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_194_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_194_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_194_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_195_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_195_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_195_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_195_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_196_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_196_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_197_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_197_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_198_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_198_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_199_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_199_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_200_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_200_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_201_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_201_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_202_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_202_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_202_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_202_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_203_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_203_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_203_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_203_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_204_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_204_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_204_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_204_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_205_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_205_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_205_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_205_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_206_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_206_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_207_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_207_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_208_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_208_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_209_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_209_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_210_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_210_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_211_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_5; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_211_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_212_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_212_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_212_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_212_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_213_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_213_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_213_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_213_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_214_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_214_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_214_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_214_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_215_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_215_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_215_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_215_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_216_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_216_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_217_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_217_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_218_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_218_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_219_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_219_io_outs_0; // @[TopModule.scala 169:11]
  wire [2:0] Multiplexer_220_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_inputs_4; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_inputs_3; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_inputs_2; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_220_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_221_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_221_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_221_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_221_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_222_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_222_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_222_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_222_io_outs_0; // @[TopModule.scala 169:11]
  wire  Multiplexer_223_io_configuration; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_223_io_inputs_1; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_223_io_inputs_0; // @[TopModule.scala 169:11]
  wire [31:0] Multiplexer_223_io_outs_0; // @[TopModule.scala 169:11]
  wire [31:0] ConstUnit_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_1_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_1_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_2_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_2_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_3_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_3_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_4_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_4_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_5_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_5_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_6_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_6_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_7_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_7_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_8_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_8_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_9_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_9_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_10_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_10_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_11_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_11_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_12_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_12_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_13_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_13_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_14_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_14_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_15_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_15_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_16_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_16_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_17_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_17_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_18_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_18_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_19_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_19_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_20_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_20_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_21_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_21_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_22_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_22_io_outs_0; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_23_io_configuration; // @[TopModule.scala 177:21]
  wire [31:0] ConstUnit_23_io_outs_0; // @[TopModule.scala 177:21]
  wire  LoadStoreUnit_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_1_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_1_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_1_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_1_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_1_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_1_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_1_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_1_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_2_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_2_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_2_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_2_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_2_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_2_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_2_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_2_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_3_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_3_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_3_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_3_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_3_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_3_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_3_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_3_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_4_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_4_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_4_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_4_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_4_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_4_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_4_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_4_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_5_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_5_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_5_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_5_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_5_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_5_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_5_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_5_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_6_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_6_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_6_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_6_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_6_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_6_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_6_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_6_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_clock; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_reset; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_configuration; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_en; // @[TopModule.scala 186:21]
  wire [3:0] LoadStoreUnit_7_io_skewing; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_streamIn_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_streamIn_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_7_io_streamIn_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_7_io_len; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_streamOut_ready; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_streamOut_valid; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_7_io_streamOut_bits; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_7_io_base; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_start; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_enqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_deqEn; // @[TopModule.scala 186:21]
  wire  LoadStoreUnit_7_io_idle; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_7_io_inputs_1; // @[TopModule.scala 186:21]
  wire [5:0] LoadStoreUnit_7_io_inputs_0; // @[TopModule.scala 186:21]
  wire [31:0] LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 186:21]
  wire  MultiIIScheduleController_16_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_16_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_16_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_16_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_16_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_16_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_16_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_17_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_17_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_17_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_17_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_17_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_17_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_17_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_18_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_18_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_18_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_18_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_18_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_18_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_18_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_19_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_19_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_19_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_19_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_19_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_19_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_19_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_20_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_20_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_20_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_20_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_20_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_20_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_20_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_21_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_21_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_21_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_21_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_21_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_21_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_21_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_22_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_22_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_22_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_22_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_22_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_22_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_22_io_skewing; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_23_clock; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_23_reset; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_23_io_en; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_0; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_1; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_2; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_3; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_4; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_5; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_6; // @[TopModule.scala 200:23]
  wire [5:0] MultiIIScheduleController_23_io_schedules_7; // @[TopModule.scala 200:23]
  wire [2:0] MultiIIScheduleController_23_io_II; // @[TopModule.scala 200:23]
  wire  MultiIIScheduleController_23_io_valid; // @[TopModule.scala 200:23]
  wire [3:0] MultiIIScheduleController_23_io_skewing; // @[TopModule.scala 200:23]
  wire  configControllers_0_clock; // @[TopModule.scala 262:34]
  wire  configControllers_0_reset; // @[TopModule.scala 262:34]
  wire  configControllers_0_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_0_io_II; // @[TopModule.scala 262:34]
  wire [35:0] configControllers_0_io_inConfig; // @[TopModule.scala 262:34]
  wire [35:0] configControllers_0_io_outConfig; // @[TopModule.scala 262:34]
  wire [35:0] Dispatch_1_io_configuration; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_1_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_1_clock; // @[TopModule.scala 262:34]
  wire  configControllers_1_reset; // @[TopModule.scala 262:34]
  wire  configControllers_1_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_1_io_II; // @[TopModule.scala 262:34]
  wire [35:0] configControllers_1_io_inConfig; // @[TopModule.scala 262:34]
  wire [35:0] configControllers_1_io_outConfig; // @[TopModule.scala 262:34]
  wire [35:0] Dispatch_2_io_configuration; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_2_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_2_clock; // @[TopModule.scala 262:34]
  wire  configControllers_2_reset; // @[TopModule.scala 262:34]
  wire  configControllers_2_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_2_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_2_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_2_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_3_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_3_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_3_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_3_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_3_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_3_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_3_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_3_clock; // @[TopModule.scala 262:34]
  wire  configControllers_3_reset; // @[TopModule.scala 262:34]
  wire  configControllers_3_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_3_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_3_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_3_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_4_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_4_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_4_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_4_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_4_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_4_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_4_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_4_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_4_clock; // @[TopModule.scala 262:34]
  wire  configControllers_4_reset; // @[TopModule.scala 262:34]
  wire  configControllers_4_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_4_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_4_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_4_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_5_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_5_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_5_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_5_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_5_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_5_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_5_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_5_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_5_clock; // @[TopModule.scala 262:34]
  wire  configControllers_5_reset; // @[TopModule.scala 262:34]
  wire  configControllers_5_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_5_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_5_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_5_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_6_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_6_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_6_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_6_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_6_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_6_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_6_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_6_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_6_clock; // @[TopModule.scala 262:34]
  wire  configControllers_6_reset; // @[TopModule.scala 262:34]
  wire  configControllers_6_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_6_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_6_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_6_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_7_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_7_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_7_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_7_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_7_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_7_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_7_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_7_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_7_clock; // @[TopModule.scala 262:34]
  wire  configControllers_7_reset; // @[TopModule.scala 262:34]
  wire  configControllers_7_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_7_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_7_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_7_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_8_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_8_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_8_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_8_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_8_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_8_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_8_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_8_clock; // @[TopModule.scala 262:34]
  wire  configControllers_8_reset; // @[TopModule.scala 262:34]
  wire  configControllers_8_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_8_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_8_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_8_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_9_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_9_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_9_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_9_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_9_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_9_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_9_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_9_clock; // @[TopModule.scala 262:34]
  wire  configControllers_9_reset; // @[TopModule.scala 262:34]
  wire  configControllers_9_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_9_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_9_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_9_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_10_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_10_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_10_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_10_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_10_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_10_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_10_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_10_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_10_clock; // @[TopModule.scala 262:34]
  wire  configControllers_10_reset; // @[TopModule.scala 262:34]
  wire  configControllers_10_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_10_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_10_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_10_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_11_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_11_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_11_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_11_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_11_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_11_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_11_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_11_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_11_clock; // @[TopModule.scala 262:34]
  wire  configControllers_11_reset; // @[TopModule.scala 262:34]
  wire  configControllers_11_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_11_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_11_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_11_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_12_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_12_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_12_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_12_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_12_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_12_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_12_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_12_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_12_clock; // @[TopModule.scala 262:34]
  wire  configControllers_12_reset; // @[TopModule.scala 262:34]
  wire  configControllers_12_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_12_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_12_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_12_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_13_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_13_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_13_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_13_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_13_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_13_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_13_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_13_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_13_clock; // @[TopModule.scala 262:34]
  wire  configControllers_13_reset; // @[TopModule.scala 262:34]
  wire  configControllers_13_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_13_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_13_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_13_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_14_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_14_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_14_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_14_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_14_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_14_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_14_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_14_clock; // @[TopModule.scala 262:34]
  wire  configControllers_14_reset; // @[TopModule.scala 262:34]
  wire  configControllers_14_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_14_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_14_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_14_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_15_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_15_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_15_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_15_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_15_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_15_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_15_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_15_clock; // @[TopModule.scala 262:34]
  wire  configControllers_15_reset; // @[TopModule.scala 262:34]
  wire  configControllers_15_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_15_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_15_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_15_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_16_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_16_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_16_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_16_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_16_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_16_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_16_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_16_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_16_clock; // @[TopModule.scala 262:34]
  wire  configControllers_16_reset; // @[TopModule.scala 262:34]
  wire  configControllers_16_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_16_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_16_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_16_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_17_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_17_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_17_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_17_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_17_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_17_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_17_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_17_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_17_clock; // @[TopModule.scala 262:34]
  wire  configControllers_17_reset; // @[TopModule.scala 262:34]
  wire  configControllers_17_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_17_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_17_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_17_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_18_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_18_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_18_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_18_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_18_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_18_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_18_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_18_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_18_clock; // @[TopModule.scala 262:34]
  wire  configControllers_18_reset; // @[TopModule.scala 262:34]
  wire  configControllers_18_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_18_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_18_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_18_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_19_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_19_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_19_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_19_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_19_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_19_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_19_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_19_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_19_clock; // @[TopModule.scala 262:34]
  wire  configControllers_19_reset; // @[TopModule.scala 262:34]
  wire  configControllers_19_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_19_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_19_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_19_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_20_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_20_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_20_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_20_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_20_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_20_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_20_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_20_clock; // @[TopModule.scala 262:34]
  wire  configControllers_20_reset; // @[TopModule.scala 262:34]
  wire  configControllers_20_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_20_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_20_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_20_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_21_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_21_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_21_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_21_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_21_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_21_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_21_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_21_clock; // @[TopModule.scala 262:34]
  wire  configControllers_21_reset; // @[TopModule.scala 262:34]
  wire  configControllers_21_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_21_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_21_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_21_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_22_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_22_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_22_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_22_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_22_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_22_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_22_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_22_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_22_clock; // @[TopModule.scala 262:34]
  wire  configControllers_22_reset; // @[TopModule.scala 262:34]
  wire  configControllers_22_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_22_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_22_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_22_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_23_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_23_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_23_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_23_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_23_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_23_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_23_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_23_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_23_clock; // @[TopModule.scala 262:34]
  wire  configControllers_23_reset; // @[TopModule.scala 262:34]
  wire  configControllers_23_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_23_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_23_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_23_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_24_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_24_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_24_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_24_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_24_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_24_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_24_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_24_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_24_clock; // @[TopModule.scala 262:34]
  wire  configControllers_24_reset; // @[TopModule.scala 262:34]
  wire  configControllers_24_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_24_io_II; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_24_io_inConfig; // @[TopModule.scala 262:34]
  wire [75:0] configControllers_24_io_outConfig; // @[TopModule.scala 262:34]
  wire [75:0] Dispatch_25_io_configuration; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_25_io_outs_17; // @[TopModule.scala 267:26]
  wire  Dispatch_25_io_outs_16; // @[TopModule.scala 267:26]
  wire  Dispatch_25_io_outs_15; // @[TopModule.scala 267:26]
  wire  Dispatch_25_io_outs_14; // @[TopModule.scala 267:26]
  wire  Dispatch_25_io_outs_13; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_12; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_11; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_10; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_9; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_25_io_outs_1; // @[TopModule.scala 267:26]
  wire [3:0] Dispatch_25_io_outs_0; // @[TopModule.scala 267:26]
  wire  configControllers_25_clock; // @[TopModule.scala 262:34]
  wire  configControllers_25_reset; // @[TopModule.scala 262:34]
  wire  configControllers_25_io_en; // @[TopModule.scala 262:34]
  wire [2:0] configControllers_25_io_II; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_25_io_inConfig; // @[TopModule.scala 262:34]
  wire [59:0] configControllers_25_io_outConfig; // @[TopModule.scala 262:34]
  wire [59:0] Dispatch_26_io_configuration; // @[TopModule.scala 267:26]
  wire  Dispatch_26_io_outs_12; // @[TopModule.scala 267:26]
  wire [31:0] Dispatch_26_io_outs_11; // @[TopModule.scala 267:26]
  wire  Dispatch_26_io_outs_10; // @[TopModule.scala 267:26]
  wire  Dispatch_26_io_outs_9; // @[TopModule.scala 267:26]
  wire  Dispatch_26_io_outs_8; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_7; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_6; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_5; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_4; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_3; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_2; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_1; // @[TopModule.scala 267:26]
  wire [2:0] Dispatch_26_io_outs_0; // @[TopModule.scala 267:26]
  wire [1767:0] topDispatch_io_configuration; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_25; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_24; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_23; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_22; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_21; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_20; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_19; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_18; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_17; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_16; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_15; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_14; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_13; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_12; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_11; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_10; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_9; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_8; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_7; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_6; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_5; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_4; // @[TopModule.scala 276:27]
  wire [75:0] topDispatch_io_outs_3; // @[TopModule.scala 276:27]
  wire [59:0] topDispatch_io_outs_2; // @[TopModule.scala 276:27]
  wire [35:0] topDispatch_io_outs_1; // @[TopModule.scala 276:27]
  wire [35:0] topDispatch_io_outs_0; // @[TopModule.scala 276:27]
  Dispatch Dispatch ( // @[TopModule.scala 122:34]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_191(Dispatch_io_outs_191),
    .io_outs_190(Dispatch_io_outs_190),
    .io_outs_189(Dispatch_io_outs_189),
    .io_outs_188(Dispatch_io_outs_188),
    .io_outs_187(Dispatch_io_outs_187),
    .io_outs_186(Dispatch_io_outs_186),
    .io_outs_185(Dispatch_io_outs_185),
    .io_outs_184(Dispatch_io_outs_184),
    .io_outs_183(Dispatch_io_outs_183),
    .io_outs_182(Dispatch_io_outs_182),
    .io_outs_181(Dispatch_io_outs_181),
    .io_outs_180(Dispatch_io_outs_180),
    .io_outs_179(Dispatch_io_outs_179),
    .io_outs_178(Dispatch_io_outs_178),
    .io_outs_177(Dispatch_io_outs_177),
    .io_outs_176(Dispatch_io_outs_176),
    .io_outs_175(Dispatch_io_outs_175),
    .io_outs_174(Dispatch_io_outs_174),
    .io_outs_173(Dispatch_io_outs_173),
    .io_outs_172(Dispatch_io_outs_172),
    .io_outs_171(Dispatch_io_outs_171),
    .io_outs_170(Dispatch_io_outs_170),
    .io_outs_169(Dispatch_io_outs_169),
    .io_outs_168(Dispatch_io_outs_168),
    .io_outs_167(Dispatch_io_outs_167),
    .io_outs_166(Dispatch_io_outs_166),
    .io_outs_165(Dispatch_io_outs_165),
    .io_outs_164(Dispatch_io_outs_164),
    .io_outs_163(Dispatch_io_outs_163),
    .io_outs_162(Dispatch_io_outs_162),
    .io_outs_161(Dispatch_io_outs_161),
    .io_outs_160(Dispatch_io_outs_160),
    .io_outs_159(Dispatch_io_outs_159),
    .io_outs_158(Dispatch_io_outs_158),
    .io_outs_157(Dispatch_io_outs_157),
    .io_outs_156(Dispatch_io_outs_156),
    .io_outs_155(Dispatch_io_outs_155),
    .io_outs_154(Dispatch_io_outs_154),
    .io_outs_153(Dispatch_io_outs_153),
    .io_outs_152(Dispatch_io_outs_152),
    .io_outs_151(Dispatch_io_outs_151),
    .io_outs_150(Dispatch_io_outs_150),
    .io_outs_149(Dispatch_io_outs_149),
    .io_outs_148(Dispatch_io_outs_148),
    .io_outs_147(Dispatch_io_outs_147),
    .io_outs_146(Dispatch_io_outs_146),
    .io_outs_145(Dispatch_io_outs_145),
    .io_outs_144(Dispatch_io_outs_144),
    .io_outs_143(Dispatch_io_outs_143),
    .io_outs_142(Dispatch_io_outs_142),
    .io_outs_141(Dispatch_io_outs_141),
    .io_outs_140(Dispatch_io_outs_140),
    .io_outs_139(Dispatch_io_outs_139),
    .io_outs_138(Dispatch_io_outs_138),
    .io_outs_137(Dispatch_io_outs_137),
    .io_outs_136(Dispatch_io_outs_136),
    .io_outs_135(Dispatch_io_outs_135),
    .io_outs_134(Dispatch_io_outs_134),
    .io_outs_133(Dispatch_io_outs_133),
    .io_outs_132(Dispatch_io_outs_132),
    .io_outs_131(Dispatch_io_outs_131),
    .io_outs_130(Dispatch_io_outs_130),
    .io_outs_129(Dispatch_io_outs_129),
    .io_outs_128(Dispatch_io_outs_128),
    .io_outs_127(Dispatch_io_outs_127),
    .io_outs_126(Dispatch_io_outs_126),
    .io_outs_125(Dispatch_io_outs_125),
    .io_outs_124(Dispatch_io_outs_124),
    .io_outs_123(Dispatch_io_outs_123),
    .io_outs_122(Dispatch_io_outs_122),
    .io_outs_121(Dispatch_io_outs_121),
    .io_outs_120(Dispatch_io_outs_120),
    .io_outs_119(Dispatch_io_outs_119),
    .io_outs_118(Dispatch_io_outs_118),
    .io_outs_117(Dispatch_io_outs_117),
    .io_outs_116(Dispatch_io_outs_116),
    .io_outs_115(Dispatch_io_outs_115),
    .io_outs_114(Dispatch_io_outs_114),
    .io_outs_113(Dispatch_io_outs_113),
    .io_outs_112(Dispatch_io_outs_112),
    .io_outs_111(Dispatch_io_outs_111),
    .io_outs_110(Dispatch_io_outs_110),
    .io_outs_109(Dispatch_io_outs_109),
    .io_outs_108(Dispatch_io_outs_108),
    .io_outs_107(Dispatch_io_outs_107),
    .io_outs_106(Dispatch_io_outs_106),
    .io_outs_105(Dispatch_io_outs_105),
    .io_outs_104(Dispatch_io_outs_104),
    .io_outs_103(Dispatch_io_outs_103),
    .io_outs_102(Dispatch_io_outs_102),
    .io_outs_101(Dispatch_io_outs_101),
    .io_outs_100(Dispatch_io_outs_100),
    .io_outs_99(Dispatch_io_outs_99),
    .io_outs_98(Dispatch_io_outs_98),
    .io_outs_97(Dispatch_io_outs_97),
    .io_outs_96(Dispatch_io_outs_96),
    .io_outs_95(Dispatch_io_outs_95),
    .io_outs_94(Dispatch_io_outs_94),
    .io_outs_93(Dispatch_io_outs_93),
    .io_outs_92(Dispatch_io_outs_92),
    .io_outs_91(Dispatch_io_outs_91),
    .io_outs_90(Dispatch_io_outs_90),
    .io_outs_89(Dispatch_io_outs_89),
    .io_outs_88(Dispatch_io_outs_88),
    .io_outs_87(Dispatch_io_outs_87),
    .io_outs_86(Dispatch_io_outs_86),
    .io_outs_85(Dispatch_io_outs_85),
    .io_outs_84(Dispatch_io_outs_84),
    .io_outs_83(Dispatch_io_outs_83),
    .io_outs_82(Dispatch_io_outs_82),
    .io_outs_81(Dispatch_io_outs_81),
    .io_outs_80(Dispatch_io_outs_80),
    .io_outs_79(Dispatch_io_outs_79),
    .io_outs_78(Dispatch_io_outs_78),
    .io_outs_77(Dispatch_io_outs_77),
    .io_outs_76(Dispatch_io_outs_76),
    .io_outs_75(Dispatch_io_outs_75),
    .io_outs_74(Dispatch_io_outs_74),
    .io_outs_73(Dispatch_io_outs_73),
    .io_outs_72(Dispatch_io_outs_72),
    .io_outs_71(Dispatch_io_outs_71),
    .io_outs_70(Dispatch_io_outs_70),
    .io_outs_69(Dispatch_io_outs_69),
    .io_outs_68(Dispatch_io_outs_68),
    .io_outs_67(Dispatch_io_outs_67),
    .io_outs_66(Dispatch_io_outs_66),
    .io_outs_65(Dispatch_io_outs_65),
    .io_outs_64(Dispatch_io_outs_64),
    .io_outs_63(Dispatch_io_outs_63),
    .io_outs_62(Dispatch_io_outs_62),
    .io_outs_61(Dispatch_io_outs_61),
    .io_outs_60(Dispatch_io_outs_60),
    .io_outs_59(Dispatch_io_outs_59),
    .io_outs_58(Dispatch_io_outs_58),
    .io_outs_57(Dispatch_io_outs_57),
    .io_outs_56(Dispatch_io_outs_56),
    .io_outs_55(Dispatch_io_outs_55),
    .io_outs_54(Dispatch_io_outs_54),
    .io_outs_53(Dispatch_io_outs_53),
    .io_outs_52(Dispatch_io_outs_52),
    .io_outs_51(Dispatch_io_outs_51),
    .io_outs_50(Dispatch_io_outs_50),
    .io_outs_49(Dispatch_io_outs_49),
    .io_outs_48(Dispatch_io_outs_48),
    .io_outs_47(Dispatch_io_outs_47),
    .io_outs_46(Dispatch_io_outs_46),
    .io_outs_45(Dispatch_io_outs_45),
    .io_outs_44(Dispatch_io_outs_44),
    .io_outs_43(Dispatch_io_outs_43),
    .io_outs_42(Dispatch_io_outs_42),
    .io_outs_41(Dispatch_io_outs_41),
    .io_outs_40(Dispatch_io_outs_40),
    .io_outs_39(Dispatch_io_outs_39),
    .io_outs_38(Dispatch_io_outs_38),
    .io_outs_37(Dispatch_io_outs_37),
    .io_outs_36(Dispatch_io_outs_36),
    .io_outs_35(Dispatch_io_outs_35),
    .io_outs_34(Dispatch_io_outs_34),
    .io_outs_33(Dispatch_io_outs_33),
    .io_outs_32(Dispatch_io_outs_32),
    .io_outs_31(Dispatch_io_outs_31),
    .io_outs_30(Dispatch_io_outs_30),
    .io_outs_29(Dispatch_io_outs_29),
    .io_outs_28(Dispatch_io_outs_28),
    .io_outs_27(Dispatch_io_outs_27),
    .io_outs_26(Dispatch_io_outs_26),
    .io_outs_25(Dispatch_io_outs_25),
    .io_outs_24(Dispatch_io_outs_24),
    .io_outs_23(Dispatch_io_outs_23),
    .io_outs_22(Dispatch_io_outs_22),
    .io_outs_21(Dispatch_io_outs_21),
    .io_outs_20(Dispatch_io_outs_20),
    .io_outs_19(Dispatch_io_outs_19),
    .io_outs_18(Dispatch_io_outs_18),
    .io_outs_17(Dispatch_io_outs_17),
    .io_outs_16(Dispatch_io_outs_16),
    .io_outs_15(Dispatch_io_outs_15),
    .io_outs_14(Dispatch_io_outs_14),
    .io_outs_13(Dispatch_io_outs_13),
    .io_outs_12(Dispatch_io_outs_12),
    .io_outs_11(Dispatch_io_outs_11),
    .io_outs_10(Dispatch_io_outs_10),
    .io_outs_9(Dispatch_io_outs_9),
    .io_outs_8(Dispatch_io_outs_8),
    .io_outs_7(Dispatch_io_outs_7),
    .io_outs_6(Dispatch_io_outs_6),
    .io_outs_5(Dispatch_io_outs_5),
    .io_outs_4(Dispatch_io_outs_4),
    .io_outs_3(Dispatch_io_outs_3),
    .io_outs_2(Dispatch_io_outs_2),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  Alu Alu ( // @[TopModule.scala 131:54]
    .clock(Alu_clock),
    .reset(Alu_reset),
    .io_en(Alu_io_en),
    .io_skewing(Alu_io_skewing),
    .io_configuration(Alu_io_configuration),
    .io_inputs_1(Alu_io_inputs_1),
    .io_inputs_0(Alu_io_inputs_0),
    .io_outs_0(Alu_io_outs_0)
  );
  Alu Alu_1 ( // @[TopModule.scala 131:54]
    .clock(Alu_1_clock),
    .reset(Alu_1_reset),
    .io_en(Alu_1_io_en),
    .io_skewing(Alu_1_io_skewing),
    .io_configuration(Alu_1_io_configuration),
    .io_inputs_1(Alu_1_io_inputs_1),
    .io_inputs_0(Alu_1_io_inputs_0),
    .io_outs_0(Alu_1_io_outs_0)
  );
  Alu Alu_2 ( // @[TopModule.scala 131:54]
    .clock(Alu_2_clock),
    .reset(Alu_2_reset),
    .io_en(Alu_2_io_en),
    .io_skewing(Alu_2_io_skewing),
    .io_configuration(Alu_2_io_configuration),
    .io_inputs_1(Alu_2_io_inputs_1),
    .io_inputs_0(Alu_2_io_inputs_0),
    .io_outs_0(Alu_2_io_outs_0)
  );
  Alu Alu_3 ( // @[TopModule.scala 131:54]
    .clock(Alu_3_clock),
    .reset(Alu_3_reset),
    .io_en(Alu_3_io_en),
    .io_skewing(Alu_3_io_skewing),
    .io_configuration(Alu_3_io_configuration),
    .io_inputs_1(Alu_3_io_inputs_1),
    .io_inputs_0(Alu_3_io_inputs_0),
    .io_outs_0(Alu_3_io_outs_0)
  );
  Alu Alu_4 ( // @[TopModule.scala 131:54]
    .clock(Alu_4_clock),
    .reset(Alu_4_reset),
    .io_en(Alu_4_io_en),
    .io_skewing(Alu_4_io_skewing),
    .io_configuration(Alu_4_io_configuration),
    .io_inputs_1(Alu_4_io_inputs_1),
    .io_inputs_0(Alu_4_io_inputs_0),
    .io_outs_0(Alu_4_io_outs_0)
  );
  Alu Alu_5 ( // @[TopModule.scala 131:54]
    .clock(Alu_5_clock),
    .reset(Alu_5_reset),
    .io_en(Alu_5_io_en),
    .io_skewing(Alu_5_io_skewing),
    .io_configuration(Alu_5_io_configuration),
    .io_inputs_1(Alu_5_io_inputs_1),
    .io_inputs_0(Alu_5_io_inputs_0),
    .io_outs_0(Alu_5_io_outs_0)
  );
  Alu Alu_6 ( // @[TopModule.scala 131:54]
    .clock(Alu_6_clock),
    .reset(Alu_6_reset),
    .io_en(Alu_6_io_en),
    .io_skewing(Alu_6_io_skewing),
    .io_configuration(Alu_6_io_configuration),
    .io_inputs_1(Alu_6_io_inputs_1),
    .io_inputs_0(Alu_6_io_inputs_0),
    .io_outs_0(Alu_6_io_outs_0)
  );
  Alu Alu_7 ( // @[TopModule.scala 131:54]
    .clock(Alu_7_clock),
    .reset(Alu_7_reset),
    .io_en(Alu_7_io_en),
    .io_skewing(Alu_7_io_skewing),
    .io_configuration(Alu_7_io_configuration),
    .io_inputs_1(Alu_7_io_inputs_1),
    .io_inputs_0(Alu_7_io_inputs_0),
    .io_outs_0(Alu_7_io_outs_0)
  );
  Alu Alu_8 ( // @[TopModule.scala 131:54]
    .clock(Alu_8_clock),
    .reset(Alu_8_reset),
    .io_en(Alu_8_io_en),
    .io_skewing(Alu_8_io_skewing),
    .io_configuration(Alu_8_io_configuration),
    .io_inputs_1(Alu_8_io_inputs_1),
    .io_inputs_0(Alu_8_io_inputs_0),
    .io_outs_0(Alu_8_io_outs_0)
  );
  Alu Alu_9 ( // @[TopModule.scala 131:54]
    .clock(Alu_9_clock),
    .reset(Alu_9_reset),
    .io_en(Alu_9_io_en),
    .io_skewing(Alu_9_io_skewing),
    .io_configuration(Alu_9_io_configuration),
    .io_inputs_1(Alu_9_io_inputs_1),
    .io_inputs_0(Alu_9_io_inputs_0),
    .io_outs_0(Alu_9_io_outs_0)
  );
  Alu Alu_10 ( // @[TopModule.scala 131:54]
    .clock(Alu_10_clock),
    .reset(Alu_10_reset),
    .io_en(Alu_10_io_en),
    .io_skewing(Alu_10_io_skewing),
    .io_configuration(Alu_10_io_configuration),
    .io_inputs_1(Alu_10_io_inputs_1),
    .io_inputs_0(Alu_10_io_inputs_0),
    .io_outs_0(Alu_10_io_outs_0)
  );
  Alu Alu_11 ( // @[TopModule.scala 131:54]
    .clock(Alu_11_clock),
    .reset(Alu_11_reset),
    .io_en(Alu_11_io_en),
    .io_skewing(Alu_11_io_skewing),
    .io_configuration(Alu_11_io_configuration),
    .io_inputs_1(Alu_11_io_inputs_1),
    .io_inputs_0(Alu_11_io_inputs_0),
    .io_outs_0(Alu_11_io_outs_0)
  );
  Alu Alu_12 ( // @[TopModule.scala 131:54]
    .clock(Alu_12_clock),
    .reset(Alu_12_reset),
    .io_en(Alu_12_io_en),
    .io_skewing(Alu_12_io_skewing),
    .io_configuration(Alu_12_io_configuration),
    .io_inputs_1(Alu_12_io_inputs_1),
    .io_inputs_0(Alu_12_io_inputs_0),
    .io_outs_0(Alu_12_io_outs_0)
  );
  Alu Alu_13 ( // @[TopModule.scala 131:54]
    .clock(Alu_13_clock),
    .reset(Alu_13_reset),
    .io_en(Alu_13_io_en),
    .io_skewing(Alu_13_io_skewing),
    .io_configuration(Alu_13_io_configuration),
    .io_inputs_1(Alu_13_io_inputs_1),
    .io_inputs_0(Alu_13_io_inputs_0),
    .io_outs_0(Alu_13_io_outs_0)
  );
  Alu Alu_14 ( // @[TopModule.scala 131:54]
    .clock(Alu_14_clock),
    .reset(Alu_14_reset),
    .io_en(Alu_14_io_en),
    .io_skewing(Alu_14_io_skewing),
    .io_configuration(Alu_14_io_configuration),
    .io_inputs_1(Alu_14_io_inputs_1),
    .io_inputs_0(Alu_14_io_inputs_0),
    .io_outs_0(Alu_14_io_outs_0)
  );
  Alu Alu_15 ( // @[TopModule.scala 131:54]
    .clock(Alu_15_clock),
    .reset(Alu_15_reset),
    .io_en(Alu_15_io_en),
    .io_skewing(Alu_15_io_skewing),
    .io_configuration(Alu_15_io_configuration),
    .io_inputs_1(Alu_15_io_inputs_1),
    .io_inputs_0(Alu_15_io_inputs_0),
    .io_outs_0(Alu_15_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_clock),
    .reset(MultiIIScheduleController_reset),
    .io_en(MultiIIScheduleController_io_en),
    .io_schedules_0(MultiIIScheduleController_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_io_schedules_7),
    .io_II(MultiIIScheduleController_io_II),
    .io_valid(MultiIIScheduleController_io_valid),
    .io_skewing(MultiIIScheduleController_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_1 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_1_clock),
    .reset(MultiIIScheduleController_1_reset),
    .io_en(MultiIIScheduleController_1_io_en),
    .io_schedules_0(MultiIIScheduleController_1_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_1_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_1_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_1_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_1_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_1_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_1_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_1_io_schedules_7),
    .io_II(MultiIIScheduleController_1_io_II),
    .io_valid(MultiIIScheduleController_1_io_valid),
    .io_skewing(MultiIIScheduleController_1_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_2 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_2_clock),
    .reset(MultiIIScheduleController_2_reset),
    .io_en(MultiIIScheduleController_2_io_en),
    .io_schedules_0(MultiIIScheduleController_2_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_2_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_2_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_2_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_2_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_2_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_2_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_2_io_schedules_7),
    .io_II(MultiIIScheduleController_2_io_II),
    .io_valid(MultiIIScheduleController_2_io_valid),
    .io_skewing(MultiIIScheduleController_2_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_3 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_3_clock),
    .reset(MultiIIScheduleController_3_reset),
    .io_en(MultiIIScheduleController_3_io_en),
    .io_schedules_0(MultiIIScheduleController_3_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_3_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_3_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_3_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_3_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_3_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_3_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_3_io_schedules_7),
    .io_II(MultiIIScheduleController_3_io_II),
    .io_valid(MultiIIScheduleController_3_io_valid),
    .io_skewing(MultiIIScheduleController_3_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_4 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_4_clock),
    .reset(MultiIIScheduleController_4_reset),
    .io_en(MultiIIScheduleController_4_io_en),
    .io_schedules_0(MultiIIScheduleController_4_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_4_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_4_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_4_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_4_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_4_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_4_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_4_io_schedules_7),
    .io_II(MultiIIScheduleController_4_io_II),
    .io_valid(MultiIIScheduleController_4_io_valid),
    .io_skewing(MultiIIScheduleController_4_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_5 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_5_clock),
    .reset(MultiIIScheduleController_5_reset),
    .io_en(MultiIIScheduleController_5_io_en),
    .io_schedules_0(MultiIIScheduleController_5_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_5_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_5_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_5_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_5_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_5_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_5_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_5_io_schedules_7),
    .io_II(MultiIIScheduleController_5_io_II),
    .io_valid(MultiIIScheduleController_5_io_valid),
    .io_skewing(MultiIIScheduleController_5_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_6 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_6_clock),
    .reset(MultiIIScheduleController_6_reset),
    .io_en(MultiIIScheduleController_6_io_en),
    .io_schedules_0(MultiIIScheduleController_6_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_6_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_6_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_6_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_6_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_6_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_6_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_6_io_schedules_7),
    .io_II(MultiIIScheduleController_6_io_II),
    .io_valid(MultiIIScheduleController_6_io_valid),
    .io_skewing(MultiIIScheduleController_6_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_7 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_7_clock),
    .reset(MultiIIScheduleController_7_reset),
    .io_en(MultiIIScheduleController_7_io_en),
    .io_schedules_0(MultiIIScheduleController_7_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_7_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_7_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_7_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_7_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_7_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_7_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_7_io_schedules_7),
    .io_II(MultiIIScheduleController_7_io_II),
    .io_valid(MultiIIScheduleController_7_io_valid),
    .io_skewing(MultiIIScheduleController_7_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_8 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_8_clock),
    .reset(MultiIIScheduleController_8_reset),
    .io_en(MultiIIScheduleController_8_io_en),
    .io_schedules_0(MultiIIScheduleController_8_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_8_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_8_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_8_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_8_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_8_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_8_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_8_io_schedules_7),
    .io_II(MultiIIScheduleController_8_io_II),
    .io_valid(MultiIIScheduleController_8_io_valid),
    .io_skewing(MultiIIScheduleController_8_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_9 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_9_clock),
    .reset(MultiIIScheduleController_9_reset),
    .io_en(MultiIIScheduleController_9_io_en),
    .io_schedules_0(MultiIIScheduleController_9_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_9_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_9_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_9_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_9_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_9_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_9_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_9_io_schedules_7),
    .io_II(MultiIIScheduleController_9_io_II),
    .io_valid(MultiIIScheduleController_9_io_valid),
    .io_skewing(MultiIIScheduleController_9_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_10 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_10_clock),
    .reset(MultiIIScheduleController_10_reset),
    .io_en(MultiIIScheduleController_10_io_en),
    .io_schedules_0(MultiIIScheduleController_10_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_10_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_10_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_10_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_10_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_10_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_10_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_10_io_schedules_7),
    .io_II(MultiIIScheduleController_10_io_II),
    .io_valid(MultiIIScheduleController_10_io_valid),
    .io_skewing(MultiIIScheduleController_10_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_11 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_11_clock),
    .reset(MultiIIScheduleController_11_reset),
    .io_en(MultiIIScheduleController_11_io_en),
    .io_schedules_0(MultiIIScheduleController_11_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_11_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_11_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_11_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_11_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_11_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_11_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_11_io_schedules_7),
    .io_II(MultiIIScheduleController_11_io_II),
    .io_valid(MultiIIScheduleController_11_io_valid),
    .io_skewing(MultiIIScheduleController_11_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_12 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_12_clock),
    .reset(MultiIIScheduleController_12_reset),
    .io_en(MultiIIScheduleController_12_io_en),
    .io_schedules_0(MultiIIScheduleController_12_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_12_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_12_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_12_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_12_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_12_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_12_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_12_io_schedules_7),
    .io_II(MultiIIScheduleController_12_io_II),
    .io_valid(MultiIIScheduleController_12_io_valid),
    .io_skewing(MultiIIScheduleController_12_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_13 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_13_clock),
    .reset(MultiIIScheduleController_13_reset),
    .io_en(MultiIIScheduleController_13_io_en),
    .io_schedules_0(MultiIIScheduleController_13_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_13_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_13_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_13_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_13_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_13_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_13_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_13_io_schedules_7),
    .io_II(MultiIIScheduleController_13_io_II),
    .io_valid(MultiIIScheduleController_13_io_valid),
    .io_skewing(MultiIIScheduleController_13_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_14 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_14_clock),
    .reset(MultiIIScheduleController_14_reset),
    .io_en(MultiIIScheduleController_14_io_en),
    .io_schedules_0(MultiIIScheduleController_14_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_14_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_14_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_14_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_14_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_14_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_14_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_14_io_schedules_7),
    .io_II(MultiIIScheduleController_14_io_II),
    .io_valid(MultiIIScheduleController_14_io_valid),
    .io_skewing(MultiIIScheduleController_14_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_15 ( // @[TopModule.scala 135:23]
    .clock(MultiIIScheduleController_15_clock),
    .reset(MultiIIScheduleController_15_reset),
    .io_en(MultiIIScheduleController_15_io_en),
    .io_schedules_0(MultiIIScheduleController_15_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_15_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_15_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_15_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_15_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_15_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_15_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_15_io_schedules_7),
    .io_II(MultiIIScheduleController_15_io_II),
    .io_valid(MultiIIScheduleController_15_io_valid),
    .io_skewing(MultiIIScheduleController_15_io_skewing)
  );
  RegisterFile RegisterFile ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_clock),
    .reset(RegisterFile_reset),
    .io_configuration(RegisterFile_io_configuration),
    .io_inputs_0(RegisterFile_io_inputs_0),
    .io_outs_0(RegisterFile_io_outs_0)
  );
  RegisterFile RegisterFile_1 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_1_clock),
    .reset(RegisterFile_1_reset),
    .io_configuration(RegisterFile_1_io_configuration),
    .io_inputs_0(RegisterFile_1_io_inputs_0),
    .io_outs_0(RegisterFile_1_io_outs_0)
  );
  RegisterFile RegisterFile_2 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_2_clock),
    .reset(RegisterFile_2_reset),
    .io_configuration(RegisterFile_2_io_configuration),
    .io_inputs_0(RegisterFile_2_io_inputs_0),
    .io_outs_0(RegisterFile_2_io_outs_0)
  );
  RegisterFile RegisterFile_3 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_3_clock),
    .reset(RegisterFile_3_reset),
    .io_configuration(RegisterFile_3_io_configuration),
    .io_inputs_0(RegisterFile_3_io_inputs_0),
    .io_outs_0(RegisterFile_3_io_outs_0)
  );
  RegisterFile RegisterFile_4 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_4_clock),
    .reset(RegisterFile_4_reset),
    .io_configuration(RegisterFile_4_io_configuration),
    .io_inputs_0(RegisterFile_4_io_inputs_0),
    .io_outs_0(RegisterFile_4_io_outs_0)
  );
  RegisterFile RegisterFile_5 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_5_clock),
    .reset(RegisterFile_5_reset),
    .io_configuration(RegisterFile_5_io_configuration),
    .io_inputs_0(RegisterFile_5_io_inputs_0),
    .io_outs_0(RegisterFile_5_io_outs_0)
  );
  RegisterFile RegisterFile_6 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_6_clock),
    .reset(RegisterFile_6_reset),
    .io_configuration(RegisterFile_6_io_configuration),
    .io_inputs_0(RegisterFile_6_io_inputs_0),
    .io_outs_0(RegisterFile_6_io_outs_0)
  );
  RegisterFile RegisterFile_7 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_7_clock),
    .reset(RegisterFile_7_reset),
    .io_configuration(RegisterFile_7_io_configuration),
    .io_inputs_0(RegisterFile_7_io_inputs_0),
    .io_outs_0(RegisterFile_7_io_outs_0)
  );
  RegisterFile RegisterFile_8 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_8_clock),
    .reset(RegisterFile_8_reset),
    .io_configuration(RegisterFile_8_io_configuration),
    .io_inputs_0(RegisterFile_8_io_inputs_0),
    .io_outs_0(RegisterFile_8_io_outs_0)
  );
  RegisterFile RegisterFile_9 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_9_clock),
    .reset(RegisterFile_9_reset),
    .io_configuration(RegisterFile_9_io_configuration),
    .io_inputs_0(RegisterFile_9_io_inputs_0),
    .io_outs_0(RegisterFile_9_io_outs_0)
  );
  RegisterFile RegisterFile_10 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_10_clock),
    .reset(RegisterFile_10_reset),
    .io_configuration(RegisterFile_10_io_configuration),
    .io_inputs_0(RegisterFile_10_io_inputs_0),
    .io_outs_0(RegisterFile_10_io_outs_0)
  );
  RegisterFile RegisterFile_11 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_11_clock),
    .reset(RegisterFile_11_reset),
    .io_configuration(RegisterFile_11_io_configuration),
    .io_inputs_0(RegisterFile_11_io_inputs_0),
    .io_outs_0(RegisterFile_11_io_outs_0)
  );
  RegisterFile RegisterFile_12 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_12_clock),
    .reset(RegisterFile_12_reset),
    .io_configuration(RegisterFile_12_io_configuration),
    .io_inputs_0(RegisterFile_12_io_inputs_0),
    .io_outs_0(RegisterFile_12_io_outs_0)
  );
  RegisterFile RegisterFile_13 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_13_clock),
    .reset(RegisterFile_13_reset),
    .io_configuration(RegisterFile_13_io_configuration),
    .io_inputs_0(RegisterFile_13_io_inputs_0),
    .io_outs_0(RegisterFile_13_io_outs_0)
  );
  RegisterFile RegisterFile_14 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_14_clock),
    .reset(RegisterFile_14_reset),
    .io_configuration(RegisterFile_14_io_configuration),
    .io_inputs_0(RegisterFile_14_io_inputs_0),
    .io_outs_0(RegisterFile_14_io_outs_0)
  );
  RegisterFile RegisterFile_15 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_15_clock),
    .reset(RegisterFile_15_reset),
    .io_configuration(RegisterFile_15_io_configuration),
    .io_inputs_0(RegisterFile_15_io_inputs_0),
    .io_outs_0(RegisterFile_15_io_outs_0)
  );
  RegisterFile RegisterFile_16 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_16_clock),
    .reset(RegisterFile_16_reset),
    .io_configuration(RegisterFile_16_io_configuration),
    .io_inputs_0(RegisterFile_16_io_inputs_0),
    .io_outs_0(RegisterFile_16_io_outs_0)
  );
  RegisterFile RegisterFile_17 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_17_clock),
    .reset(RegisterFile_17_reset),
    .io_configuration(RegisterFile_17_io_configuration),
    .io_inputs_0(RegisterFile_17_io_inputs_0),
    .io_outs_0(RegisterFile_17_io_outs_0)
  );
  RegisterFile RegisterFile_18 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_18_clock),
    .reset(RegisterFile_18_reset),
    .io_configuration(RegisterFile_18_io_configuration),
    .io_inputs_0(RegisterFile_18_io_inputs_0),
    .io_outs_0(RegisterFile_18_io_outs_0)
  );
  RegisterFile RegisterFile_19 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_19_clock),
    .reset(RegisterFile_19_reset),
    .io_configuration(RegisterFile_19_io_configuration),
    .io_inputs_0(RegisterFile_19_io_inputs_0),
    .io_outs_0(RegisterFile_19_io_outs_0)
  );
  RegisterFile RegisterFile_20 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_20_clock),
    .reset(RegisterFile_20_reset),
    .io_configuration(RegisterFile_20_io_configuration),
    .io_inputs_0(RegisterFile_20_io_inputs_0),
    .io_outs_0(RegisterFile_20_io_outs_0)
  );
  RegisterFile RegisterFile_21 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_21_clock),
    .reset(RegisterFile_21_reset),
    .io_configuration(RegisterFile_21_io_configuration),
    .io_inputs_0(RegisterFile_21_io_inputs_0),
    .io_outs_0(RegisterFile_21_io_outs_0)
  );
  RegisterFile RegisterFile_22 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_22_clock),
    .reset(RegisterFile_22_reset),
    .io_configuration(RegisterFile_22_io_configuration),
    .io_inputs_0(RegisterFile_22_io_inputs_0),
    .io_outs_0(RegisterFile_22_io_outs_0)
  );
  RegisterFile RegisterFile_23 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_23_clock),
    .reset(RegisterFile_23_reset),
    .io_configuration(RegisterFile_23_io_configuration),
    .io_inputs_0(RegisterFile_23_io_inputs_0),
    .io_outs_0(RegisterFile_23_io_outs_0)
  );
  RegisterFile RegisterFile_24 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_24_clock),
    .reset(RegisterFile_24_reset),
    .io_configuration(RegisterFile_24_io_configuration),
    .io_inputs_0(RegisterFile_24_io_inputs_0),
    .io_outs_0(RegisterFile_24_io_outs_0)
  );
  RegisterFile RegisterFile_25 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_25_clock),
    .reset(RegisterFile_25_reset),
    .io_configuration(RegisterFile_25_io_configuration),
    .io_inputs_0(RegisterFile_25_io_inputs_0),
    .io_outs_0(RegisterFile_25_io_outs_0)
  );
  RegisterFile RegisterFile_26 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_26_clock),
    .reset(RegisterFile_26_reset),
    .io_configuration(RegisterFile_26_io_configuration),
    .io_inputs_0(RegisterFile_26_io_inputs_0),
    .io_outs_0(RegisterFile_26_io_outs_0)
  );
  RegisterFile RegisterFile_27 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_27_clock),
    .reset(RegisterFile_27_reset),
    .io_configuration(RegisterFile_27_io_configuration),
    .io_inputs_0(RegisterFile_27_io_inputs_0),
    .io_outs_0(RegisterFile_27_io_outs_0)
  );
  RegisterFile RegisterFile_28 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_28_clock),
    .reset(RegisterFile_28_reset),
    .io_configuration(RegisterFile_28_io_configuration),
    .io_inputs_0(RegisterFile_28_io_inputs_0),
    .io_outs_0(RegisterFile_28_io_outs_0)
  );
  RegisterFile RegisterFile_29 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_29_clock),
    .reset(RegisterFile_29_reset),
    .io_configuration(RegisterFile_29_io_configuration),
    .io_inputs_0(RegisterFile_29_io_inputs_0),
    .io_outs_0(RegisterFile_29_io_outs_0)
  );
  RegisterFile RegisterFile_30 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_30_clock),
    .reset(RegisterFile_30_reset),
    .io_configuration(RegisterFile_30_io_configuration),
    .io_inputs_0(RegisterFile_30_io_inputs_0),
    .io_outs_0(RegisterFile_30_io_outs_0)
  );
  RegisterFile RegisterFile_31 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_31_clock),
    .reset(RegisterFile_31_reset),
    .io_configuration(RegisterFile_31_io_configuration),
    .io_inputs_0(RegisterFile_31_io_inputs_0),
    .io_outs_0(RegisterFile_31_io_outs_0)
  );
  RegisterFile RegisterFile_32 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_32_clock),
    .reset(RegisterFile_32_reset),
    .io_configuration(RegisterFile_32_io_configuration),
    .io_inputs_0(RegisterFile_32_io_inputs_0),
    .io_outs_0(RegisterFile_32_io_outs_0)
  );
  RegisterFile RegisterFile_33 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_33_clock),
    .reset(RegisterFile_33_reset),
    .io_configuration(RegisterFile_33_io_configuration),
    .io_inputs_0(RegisterFile_33_io_inputs_0),
    .io_outs_0(RegisterFile_33_io_outs_0)
  );
  RegisterFile RegisterFile_34 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_34_clock),
    .reset(RegisterFile_34_reset),
    .io_configuration(RegisterFile_34_io_configuration),
    .io_inputs_0(RegisterFile_34_io_inputs_0),
    .io_outs_0(RegisterFile_34_io_outs_0)
  );
  RegisterFile RegisterFile_35 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_35_clock),
    .reset(RegisterFile_35_reset),
    .io_configuration(RegisterFile_35_io_configuration),
    .io_inputs_0(RegisterFile_35_io_inputs_0),
    .io_outs_0(RegisterFile_35_io_outs_0)
  );
  RegisterFile RegisterFile_36 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_36_clock),
    .reset(RegisterFile_36_reset),
    .io_configuration(RegisterFile_36_io_configuration),
    .io_inputs_0(RegisterFile_36_io_inputs_0),
    .io_outs_0(RegisterFile_36_io_outs_0)
  );
  RegisterFile RegisterFile_37 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_37_clock),
    .reset(RegisterFile_37_reset),
    .io_configuration(RegisterFile_37_io_configuration),
    .io_inputs_0(RegisterFile_37_io_inputs_0),
    .io_outs_0(RegisterFile_37_io_outs_0)
  );
  RegisterFile RegisterFile_38 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_38_clock),
    .reset(RegisterFile_38_reset),
    .io_configuration(RegisterFile_38_io_configuration),
    .io_inputs_0(RegisterFile_38_io_inputs_0),
    .io_outs_0(RegisterFile_38_io_outs_0)
  );
  RegisterFile RegisterFile_39 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_39_clock),
    .reset(RegisterFile_39_reset),
    .io_configuration(RegisterFile_39_io_configuration),
    .io_inputs_0(RegisterFile_39_io_inputs_0),
    .io_outs_0(RegisterFile_39_io_outs_0)
  );
  RegisterFile RegisterFile_40 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_40_clock),
    .reset(RegisterFile_40_reset),
    .io_configuration(RegisterFile_40_io_configuration),
    .io_inputs_0(RegisterFile_40_io_inputs_0),
    .io_outs_0(RegisterFile_40_io_outs_0)
  );
  RegisterFile RegisterFile_41 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_41_clock),
    .reset(RegisterFile_41_reset),
    .io_configuration(RegisterFile_41_io_configuration),
    .io_inputs_0(RegisterFile_41_io_inputs_0),
    .io_outs_0(RegisterFile_41_io_outs_0)
  );
  RegisterFile RegisterFile_42 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_42_clock),
    .reset(RegisterFile_42_reset),
    .io_configuration(RegisterFile_42_io_configuration),
    .io_inputs_0(RegisterFile_42_io_inputs_0),
    .io_outs_0(RegisterFile_42_io_outs_0)
  );
  RegisterFile RegisterFile_43 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_43_clock),
    .reset(RegisterFile_43_reset),
    .io_configuration(RegisterFile_43_io_configuration),
    .io_inputs_0(RegisterFile_43_io_inputs_0),
    .io_outs_0(RegisterFile_43_io_outs_0)
  );
  RegisterFile RegisterFile_44 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_44_clock),
    .reset(RegisterFile_44_reset),
    .io_configuration(RegisterFile_44_io_configuration),
    .io_inputs_0(RegisterFile_44_io_inputs_0),
    .io_outs_0(RegisterFile_44_io_outs_0)
  );
  RegisterFile RegisterFile_45 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_45_clock),
    .reset(RegisterFile_45_reset),
    .io_configuration(RegisterFile_45_io_configuration),
    .io_inputs_0(RegisterFile_45_io_inputs_0),
    .io_outs_0(RegisterFile_45_io_outs_0)
  );
  RegisterFile RegisterFile_46 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_46_clock),
    .reset(RegisterFile_46_reset),
    .io_configuration(RegisterFile_46_io_configuration),
    .io_inputs_0(RegisterFile_46_io_inputs_0),
    .io_outs_0(RegisterFile_46_io_outs_0)
  );
  RegisterFile RegisterFile_47 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_47_clock),
    .reset(RegisterFile_47_reset),
    .io_configuration(RegisterFile_47_io_configuration),
    .io_inputs_0(RegisterFile_47_io_inputs_0),
    .io_outs_0(RegisterFile_47_io_outs_0)
  );
  RegisterFile RegisterFile_48 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_48_clock),
    .reset(RegisterFile_48_reset),
    .io_configuration(RegisterFile_48_io_configuration),
    .io_inputs_0(RegisterFile_48_io_inputs_0),
    .io_outs_0(RegisterFile_48_io_outs_0)
  );
  RegisterFile RegisterFile_49 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_49_clock),
    .reset(RegisterFile_49_reset),
    .io_configuration(RegisterFile_49_io_configuration),
    .io_inputs_0(RegisterFile_49_io_inputs_0),
    .io_outs_0(RegisterFile_49_io_outs_0)
  );
  RegisterFile RegisterFile_50 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_50_clock),
    .reset(RegisterFile_50_reset),
    .io_configuration(RegisterFile_50_io_configuration),
    .io_inputs_0(RegisterFile_50_io_inputs_0),
    .io_outs_0(RegisterFile_50_io_outs_0)
  );
  RegisterFile RegisterFile_51 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_51_clock),
    .reset(RegisterFile_51_reset),
    .io_configuration(RegisterFile_51_io_configuration),
    .io_inputs_0(RegisterFile_51_io_inputs_0),
    .io_outs_0(RegisterFile_51_io_outs_0)
  );
  RegisterFile RegisterFile_52 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_52_clock),
    .reset(RegisterFile_52_reset),
    .io_configuration(RegisterFile_52_io_configuration),
    .io_inputs_0(RegisterFile_52_io_inputs_0),
    .io_outs_0(RegisterFile_52_io_outs_0)
  );
  RegisterFile RegisterFile_53 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_53_clock),
    .reset(RegisterFile_53_reset),
    .io_configuration(RegisterFile_53_io_configuration),
    .io_inputs_0(RegisterFile_53_io_inputs_0),
    .io_outs_0(RegisterFile_53_io_outs_0)
  );
  RegisterFile RegisterFile_54 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_54_clock),
    .reset(RegisterFile_54_reset),
    .io_configuration(RegisterFile_54_io_configuration),
    .io_inputs_0(RegisterFile_54_io_inputs_0),
    .io_outs_0(RegisterFile_54_io_outs_0)
  );
  RegisterFile RegisterFile_55 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_55_clock),
    .reset(RegisterFile_55_reset),
    .io_configuration(RegisterFile_55_io_configuration),
    .io_inputs_0(RegisterFile_55_io_inputs_0),
    .io_outs_0(RegisterFile_55_io_outs_0)
  );
  RegisterFile RegisterFile_56 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_56_clock),
    .reset(RegisterFile_56_reset),
    .io_configuration(RegisterFile_56_io_configuration),
    .io_inputs_0(RegisterFile_56_io_inputs_0),
    .io_outs_0(RegisterFile_56_io_outs_0)
  );
  RegisterFile RegisterFile_57 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_57_clock),
    .reset(RegisterFile_57_reset),
    .io_configuration(RegisterFile_57_io_configuration),
    .io_inputs_0(RegisterFile_57_io_inputs_0),
    .io_outs_0(RegisterFile_57_io_outs_0)
  );
  RegisterFile RegisterFile_58 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_58_clock),
    .reset(RegisterFile_58_reset),
    .io_configuration(RegisterFile_58_io_configuration),
    .io_inputs_0(RegisterFile_58_io_inputs_0),
    .io_outs_0(RegisterFile_58_io_outs_0)
  );
  RegisterFile RegisterFile_59 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_59_clock),
    .reset(RegisterFile_59_reset),
    .io_configuration(RegisterFile_59_io_configuration),
    .io_inputs_0(RegisterFile_59_io_inputs_0),
    .io_outs_0(RegisterFile_59_io_outs_0)
  );
  RegisterFile RegisterFile_60 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_60_clock),
    .reset(RegisterFile_60_reset),
    .io_configuration(RegisterFile_60_io_configuration),
    .io_inputs_0(RegisterFile_60_io_inputs_0),
    .io_outs_0(RegisterFile_60_io_outs_0)
  );
  RegisterFile RegisterFile_61 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_61_clock),
    .reset(RegisterFile_61_reset),
    .io_configuration(RegisterFile_61_io_configuration),
    .io_inputs_0(RegisterFile_61_io_inputs_0),
    .io_outs_0(RegisterFile_61_io_outs_0)
  );
  RegisterFile RegisterFile_62 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_62_clock),
    .reset(RegisterFile_62_reset),
    .io_configuration(RegisterFile_62_io_configuration),
    .io_inputs_0(RegisterFile_62_io_inputs_0),
    .io_outs_0(RegisterFile_62_io_outs_0)
  );
  RegisterFile RegisterFile_63 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_63_clock),
    .reset(RegisterFile_63_reset),
    .io_configuration(RegisterFile_63_io_configuration),
    .io_inputs_0(RegisterFile_63_io_inputs_0),
    .io_outs_0(RegisterFile_63_io_outs_0)
  );
  RegisterFile RegisterFile_64 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_64_clock),
    .reset(RegisterFile_64_reset),
    .io_configuration(RegisterFile_64_io_configuration),
    .io_inputs_0(RegisterFile_64_io_inputs_0),
    .io_outs_0(RegisterFile_64_io_outs_0)
  );
  RegisterFile RegisterFile_65 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_65_clock),
    .reset(RegisterFile_65_reset),
    .io_configuration(RegisterFile_65_io_configuration),
    .io_inputs_0(RegisterFile_65_io_inputs_0),
    .io_outs_0(RegisterFile_65_io_outs_0)
  );
  RegisterFile RegisterFile_66 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_66_clock),
    .reset(RegisterFile_66_reset),
    .io_configuration(RegisterFile_66_io_configuration),
    .io_inputs_0(RegisterFile_66_io_inputs_0),
    .io_outs_0(RegisterFile_66_io_outs_0)
  );
  RegisterFile RegisterFile_67 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_67_clock),
    .reset(RegisterFile_67_reset),
    .io_configuration(RegisterFile_67_io_configuration),
    .io_inputs_0(RegisterFile_67_io_inputs_0),
    .io_outs_0(RegisterFile_67_io_outs_0)
  );
  RegisterFile RegisterFile_68 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_68_clock),
    .reset(RegisterFile_68_reset),
    .io_configuration(RegisterFile_68_io_configuration),
    .io_inputs_0(RegisterFile_68_io_inputs_0),
    .io_outs_0(RegisterFile_68_io_outs_0)
  );
  RegisterFile RegisterFile_69 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_69_clock),
    .reset(RegisterFile_69_reset),
    .io_configuration(RegisterFile_69_io_configuration),
    .io_inputs_0(RegisterFile_69_io_inputs_0),
    .io_outs_0(RegisterFile_69_io_outs_0)
  );
  RegisterFile RegisterFile_70 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_70_clock),
    .reset(RegisterFile_70_reset),
    .io_configuration(RegisterFile_70_io_configuration),
    .io_inputs_0(RegisterFile_70_io_inputs_0),
    .io_outs_0(RegisterFile_70_io_outs_0)
  );
  RegisterFile RegisterFile_71 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_71_clock),
    .reset(RegisterFile_71_reset),
    .io_configuration(RegisterFile_71_io_configuration),
    .io_inputs_0(RegisterFile_71_io_inputs_0),
    .io_outs_0(RegisterFile_71_io_outs_0)
  );
  RegisterFile RegisterFile_72 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_72_clock),
    .reset(RegisterFile_72_reset),
    .io_configuration(RegisterFile_72_io_configuration),
    .io_inputs_0(RegisterFile_72_io_inputs_0),
    .io_outs_0(RegisterFile_72_io_outs_0)
  );
  RegisterFile RegisterFile_73 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_73_clock),
    .reset(RegisterFile_73_reset),
    .io_configuration(RegisterFile_73_io_configuration),
    .io_inputs_0(RegisterFile_73_io_inputs_0),
    .io_outs_0(RegisterFile_73_io_outs_0)
  );
  RegisterFile RegisterFile_74 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_74_clock),
    .reset(RegisterFile_74_reset),
    .io_configuration(RegisterFile_74_io_configuration),
    .io_inputs_0(RegisterFile_74_io_inputs_0),
    .io_outs_0(RegisterFile_74_io_outs_0)
  );
  RegisterFile RegisterFile_75 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_75_clock),
    .reset(RegisterFile_75_reset),
    .io_configuration(RegisterFile_75_io_configuration),
    .io_inputs_0(RegisterFile_75_io_inputs_0),
    .io_outs_0(RegisterFile_75_io_outs_0)
  );
  RegisterFile RegisterFile_76 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_76_clock),
    .reset(RegisterFile_76_reset),
    .io_configuration(RegisterFile_76_io_configuration),
    .io_inputs_0(RegisterFile_76_io_inputs_0),
    .io_outs_0(RegisterFile_76_io_outs_0)
  );
  RegisterFile RegisterFile_77 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_77_clock),
    .reset(RegisterFile_77_reset),
    .io_configuration(RegisterFile_77_io_configuration),
    .io_inputs_0(RegisterFile_77_io_inputs_0),
    .io_outs_0(RegisterFile_77_io_outs_0)
  );
  RegisterFile RegisterFile_78 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_78_clock),
    .reset(RegisterFile_78_reset),
    .io_configuration(RegisterFile_78_io_configuration),
    .io_inputs_0(RegisterFile_78_io_inputs_0),
    .io_outs_0(RegisterFile_78_io_outs_0)
  );
  RegisterFile RegisterFile_79 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_79_clock),
    .reset(RegisterFile_79_reset),
    .io_configuration(RegisterFile_79_io_configuration),
    .io_inputs_0(RegisterFile_79_io_inputs_0),
    .io_outs_0(RegisterFile_79_io_outs_0)
  );
  RegisterFile RegisterFile_80 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_80_clock),
    .reset(RegisterFile_80_reset),
    .io_configuration(RegisterFile_80_io_configuration),
    .io_inputs_0(RegisterFile_80_io_inputs_0),
    .io_outs_0(RegisterFile_80_io_outs_0)
  );
  RegisterFile RegisterFile_81 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_81_clock),
    .reset(RegisterFile_81_reset),
    .io_configuration(RegisterFile_81_io_configuration),
    .io_inputs_0(RegisterFile_81_io_inputs_0),
    .io_outs_0(RegisterFile_81_io_outs_0)
  );
  RegisterFile RegisterFile_82 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_82_clock),
    .reset(RegisterFile_82_reset),
    .io_configuration(RegisterFile_82_io_configuration),
    .io_inputs_0(RegisterFile_82_io_inputs_0),
    .io_outs_0(RegisterFile_82_io_outs_0)
  );
  RegisterFile RegisterFile_83 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_83_clock),
    .reset(RegisterFile_83_reset),
    .io_configuration(RegisterFile_83_io_configuration),
    .io_inputs_0(RegisterFile_83_io_inputs_0),
    .io_outs_0(RegisterFile_83_io_outs_0)
  );
  RegisterFile RegisterFile_84 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_84_clock),
    .reset(RegisterFile_84_reset),
    .io_configuration(RegisterFile_84_io_configuration),
    .io_inputs_0(RegisterFile_84_io_inputs_0),
    .io_outs_0(RegisterFile_84_io_outs_0)
  );
  RegisterFile RegisterFile_85 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_85_clock),
    .reset(RegisterFile_85_reset),
    .io_configuration(RegisterFile_85_io_configuration),
    .io_inputs_0(RegisterFile_85_io_inputs_0),
    .io_outs_0(RegisterFile_85_io_outs_0)
  );
  RegisterFile RegisterFile_86 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_86_clock),
    .reset(RegisterFile_86_reset),
    .io_configuration(RegisterFile_86_io_configuration),
    .io_inputs_0(RegisterFile_86_io_inputs_0),
    .io_outs_0(RegisterFile_86_io_outs_0)
  );
  RegisterFile RegisterFile_87 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_87_clock),
    .reset(RegisterFile_87_reset),
    .io_configuration(RegisterFile_87_io_configuration),
    .io_inputs_0(RegisterFile_87_io_inputs_0),
    .io_outs_0(RegisterFile_87_io_outs_0)
  );
  RegisterFile RegisterFile_88 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_88_clock),
    .reset(RegisterFile_88_reset),
    .io_configuration(RegisterFile_88_io_configuration),
    .io_inputs_0(RegisterFile_88_io_inputs_0),
    .io_outs_0(RegisterFile_88_io_outs_0)
  );
  RegisterFile RegisterFile_89 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_89_clock),
    .reset(RegisterFile_89_reset),
    .io_configuration(RegisterFile_89_io_configuration),
    .io_inputs_0(RegisterFile_89_io_inputs_0),
    .io_outs_0(RegisterFile_89_io_outs_0)
  );
  RegisterFile RegisterFile_90 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_90_clock),
    .reset(RegisterFile_90_reset),
    .io_configuration(RegisterFile_90_io_configuration),
    .io_inputs_0(RegisterFile_90_io_inputs_0),
    .io_outs_0(RegisterFile_90_io_outs_0)
  );
  RegisterFile RegisterFile_91 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_91_clock),
    .reset(RegisterFile_91_reset),
    .io_configuration(RegisterFile_91_io_configuration),
    .io_inputs_0(RegisterFile_91_io_inputs_0),
    .io_outs_0(RegisterFile_91_io_outs_0)
  );
  RegisterFile RegisterFile_92 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_92_clock),
    .reset(RegisterFile_92_reset),
    .io_configuration(RegisterFile_92_io_configuration),
    .io_inputs_0(RegisterFile_92_io_inputs_0),
    .io_outs_0(RegisterFile_92_io_outs_0)
  );
  RegisterFile RegisterFile_93 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_93_clock),
    .reset(RegisterFile_93_reset),
    .io_configuration(RegisterFile_93_io_configuration),
    .io_inputs_0(RegisterFile_93_io_inputs_0),
    .io_outs_0(RegisterFile_93_io_outs_0)
  );
  RegisterFile RegisterFile_94 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_94_clock),
    .reset(RegisterFile_94_reset),
    .io_configuration(RegisterFile_94_io_configuration),
    .io_inputs_0(RegisterFile_94_io_inputs_0),
    .io_outs_0(RegisterFile_94_io_outs_0)
  );
  RegisterFile RegisterFile_95 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_95_clock),
    .reset(RegisterFile_95_reset),
    .io_configuration(RegisterFile_95_io_configuration),
    .io_inputs_0(RegisterFile_95_io_inputs_0),
    .io_outs_0(RegisterFile_95_io_outs_0)
  );
  RegisterFile RegisterFile_96 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_96_clock),
    .reset(RegisterFile_96_reset),
    .io_configuration(RegisterFile_96_io_configuration),
    .io_inputs_0(RegisterFile_96_io_inputs_0),
    .io_outs_0(RegisterFile_96_io_outs_0)
  );
  RegisterFile RegisterFile_97 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_97_clock),
    .reset(RegisterFile_97_reset),
    .io_configuration(RegisterFile_97_io_configuration),
    .io_inputs_0(RegisterFile_97_io_inputs_0),
    .io_outs_0(RegisterFile_97_io_outs_0)
  );
  RegisterFile RegisterFile_98 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_98_clock),
    .reset(RegisterFile_98_reset),
    .io_configuration(RegisterFile_98_io_configuration),
    .io_inputs_0(RegisterFile_98_io_inputs_0),
    .io_outs_0(RegisterFile_98_io_outs_0)
  );
  RegisterFile RegisterFile_99 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_99_clock),
    .reset(RegisterFile_99_reset),
    .io_configuration(RegisterFile_99_io_configuration),
    .io_inputs_0(RegisterFile_99_io_inputs_0),
    .io_outs_0(RegisterFile_99_io_outs_0)
  );
  RegisterFile RegisterFile_100 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_100_clock),
    .reset(RegisterFile_100_reset),
    .io_configuration(RegisterFile_100_io_configuration),
    .io_inputs_0(RegisterFile_100_io_inputs_0),
    .io_outs_0(RegisterFile_100_io_outs_0)
  );
  RegisterFile RegisterFile_101 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_101_clock),
    .reset(RegisterFile_101_reset),
    .io_configuration(RegisterFile_101_io_configuration),
    .io_inputs_0(RegisterFile_101_io_inputs_0),
    .io_outs_0(RegisterFile_101_io_outs_0)
  );
  RegisterFile RegisterFile_102 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_102_clock),
    .reset(RegisterFile_102_reset),
    .io_configuration(RegisterFile_102_io_configuration),
    .io_inputs_0(RegisterFile_102_io_inputs_0),
    .io_outs_0(RegisterFile_102_io_outs_0)
  );
  RegisterFile RegisterFile_103 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_103_clock),
    .reset(RegisterFile_103_reset),
    .io_configuration(RegisterFile_103_io_configuration),
    .io_inputs_0(RegisterFile_103_io_inputs_0),
    .io_outs_0(RegisterFile_103_io_outs_0)
  );
  RegisterFile RegisterFile_104 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_104_clock),
    .reset(RegisterFile_104_reset),
    .io_configuration(RegisterFile_104_io_configuration),
    .io_inputs_0(RegisterFile_104_io_inputs_0),
    .io_outs_0(RegisterFile_104_io_outs_0)
  );
  RegisterFile RegisterFile_105 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_105_clock),
    .reset(RegisterFile_105_reset),
    .io_configuration(RegisterFile_105_io_configuration),
    .io_inputs_0(RegisterFile_105_io_inputs_0),
    .io_outs_0(RegisterFile_105_io_outs_0)
  );
  RegisterFile RegisterFile_106 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_106_clock),
    .reset(RegisterFile_106_reset),
    .io_configuration(RegisterFile_106_io_configuration),
    .io_inputs_0(RegisterFile_106_io_inputs_0),
    .io_outs_0(RegisterFile_106_io_outs_0)
  );
  RegisterFile RegisterFile_107 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_107_clock),
    .reset(RegisterFile_107_reset),
    .io_configuration(RegisterFile_107_io_configuration),
    .io_inputs_0(RegisterFile_107_io_inputs_0),
    .io_outs_0(RegisterFile_107_io_outs_0)
  );
  RegisterFile RegisterFile_108 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_108_clock),
    .reset(RegisterFile_108_reset),
    .io_configuration(RegisterFile_108_io_configuration),
    .io_inputs_0(RegisterFile_108_io_inputs_0),
    .io_outs_0(RegisterFile_108_io_outs_0)
  );
  RegisterFile RegisterFile_109 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_109_clock),
    .reset(RegisterFile_109_reset),
    .io_configuration(RegisterFile_109_io_configuration),
    .io_inputs_0(RegisterFile_109_io_inputs_0),
    .io_outs_0(RegisterFile_109_io_outs_0)
  );
  RegisterFile RegisterFile_110 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_110_clock),
    .reset(RegisterFile_110_reset),
    .io_configuration(RegisterFile_110_io_configuration),
    .io_inputs_0(RegisterFile_110_io_inputs_0),
    .io_outs_0(RegisterFile_110_io_outs_0)
  );
  RegisterFile RegisterFile_111 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_111_clock),
    .reset(RegisterFile_111_reset),
    .io_configuration(RegisterFile_111_io_configuration),
    .io_inputs_0(RegisterFile_111_io_inputs_0),
    .io_outs_0(RegisterFile_111_io_outs_0)
  );
  RegisterFile RegisterFile_112 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_112_clock),
    .reset(RegisterFile_112_reset),
    .io_configuration(RegisterFile_112_io_configuration),
    .io_inputs_0(RegisterFile_112_io_inputs_0),
    .io_outs_0(RegisterFile_112_io_outs_0)
  );
  RegisterFile RegisterFile_113 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_113_clock),
    .reset(RegisterFile_113_reset),
    .io_configuration(RegisterFile_113_io_configuration),
    .io_inputs_0(RegisterFile_113_io_inputs_0),
    .io_outs_0(RegisterFile_113_io_outs_0)
  );
  RegisterFile RegisterFile_114 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_114_clock),
    .reset(RegisterFile_114_reset),
    .io_configuration(RegisterFile_114_io_configuration),
    .io_inputs_0(RegisterFile_114_io_inputs_0),
    .io_outs_0(RegisterFile_114_io_outs_0)
  );
  RegisterFile RegisterFile_115 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_115_clock),
    .reset(RegisterFile_115_reset),
    .io_configuration(RegisterFile_115_io_configuration),
    .io_inputs_0(RegisterFile_115_io_inputs_0),
    .io_outs_0(RegisterFile_115_io_outs_0)
  );
  RegisterFile RegisterFile_116 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_116_clock),
    .reset(RegisterFile_116_reset),
    .io_configuration(RegisterFile_116_io_configuration),
    .io_inputs_0(RegisterFile_116_io_inputs_0),
    .io_outs_0(RegisterFile_116_io_outs_0)
  );
  RegisterFile RegisterFile_117 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_117_clock),
    .reset(RegisterFile_117_reset),
    .io_configuration(RegisterFile_117_io_configuration),
    .io_inputs_0(RegisterFile_117_io_inputs_0),
    .io_outs_0(RegisterFile_117_io_outs_0)
  );
  RegisterFile RegisterFile_118 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_118_clock),
    .reset(RegisterFile_118_reset),
    .io_configuration(RegisterFile_118_io_configuration),
    .io_inputs_0(RegisterFile_118_io_inputs_0),
    .io_outs_0(RegisterFile_118_io_outs_0)
  );
  RegisterFile RegisterFile_119 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_119_clock),
    .reset(RegisterFile_119_reset),
    .io_configuration(RegisterFile_119_io_configuration),
    .io_inputs_0(RegisterFile_119_io_inputs_0),
    .io_outs_0(RegisterFile_119_io_outs_0)
  );
  RegisterFile RegisterFile_120 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_120_clock),
    .reset(RegisterFile_120_reset),
    .io_configuration(RegisterFile_120_io_configuration),
    .io_inputs_0(RegisterFile_120_io_inputs_0),
    .io_outs_0(RegisterFile_120_io_outs_0)
  );
  RegisterFile RegisterFile_121 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_121_clock),
    .reset(RegisterFile_121_reset),
    .io_configuration(RegisterFile_121_io_configuration),
    .io_inputs_0(RegisterFile_121_io_inputs_0),
    .io_outs_0(RegisterFile_121_io_outs_0)
  );
  RegisterFile RegisterFile_122 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_122_clock),
    .reset(RegisterFile_122_reset),
    .io_configuration(RegisterFile_122_io_configuration),
    .io_inputs_0(RegisterFile_122_io_inputs_0),
    .io_outs_0(RegisterFile_122_io_outs_0)
  );
  RegisterFile RegisterFile_123 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_123_clock),
    .reset(RegisterFile_123_reset),
    .io_configuration(RegisterFile_123_io_configuration),
    .io_inputs_0(RegisterFile_123_io_inputs_0),
    .io_outs_0(RegisterFile_123_io_outs_0)
  );
  RegisterFile RegisterFile_124 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_124_clock),
    .reset(RegisterFile_124_reset),
    .io_configuration(RegisterFile_124_io_configuration),
    .io_inputs_0(RegisterFile_124_io_inputs_0),
    .io_outs_0(RegisterFile_124_io_outs_0)
  );
  RegisterFile RegisterFile_125 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_125_clock),
    .reset(RegisterFile_125_reset),
    .io_configuration(RegisterFile_125_io_configuration),
    .io_inputs_0(RegisterFile_125_io_inputs_0),
    .io_outs_0(RegisterFile_125_io_outs_0)
  );
  RegisterFile RegisterFile_126 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_126_clock),
    .reset(RegisterFile_126_reset),
    .io_configuration(RegisterFile_126_io_configuration),
    .io_inputs_0(RegisterFile_126_io_inputs_0),
    .io_outs_0(RegisterFile_126_io_outs_0)
  );
  RegisterFile RegisterFile_127 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_127_clock),
    .reset(RegisterFile_127_reset),
    .io_configuration(RegisterFile_127_io_configuration),
    .io_inputs_0(RegisterFile_127_io_inputs_0),
    .io_outs_0(RegisterFile_127_io_outs_0)
  );
  RegisterFile RegisterFile_128 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_128_clock),
    .reset(RegisterFile_128_reset),
    .io_configuration(RegisterFile_128_io_configuration),
    .io_inputs_0(RegisterFile_128_io_inputs_0),
    .io_outs_0(RegisterFile_128_io_outs_0)
  );
  RegisterFile RegisterFile_129 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_129_clock),
    .reset(RegisterFile_129_reset),
    .io_configuration(RegisterFile_129_io_configuration),
    .io_inputs_0(RegisterFile_129_io_inputs_0),
    .io_outs_0(RegisterFile_129_io_outs_0)
  );
  RegisterFile RegisterFile_130 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_130_clock),
    .reset(RegisterFile_130_reset),
    .io_configuration(RegisterFile_130_io_configuration),
    .io_inputs_0(RegisterFile_130_io_inputs_0),
    .io_outs_0(RegisterFile_130_io_outs_0)
  );
  RegisterFile RegisterFile_131 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_131_clock),
    .reset(RegisterFile_131_reset),
    .io_configuration(RegisterFile_131_io_configuration),
    .io_inputs_0(RegisterFile_131_io_inputs_0),
    .io_outs_0(RegisterFile_131_io_outs_0)
  );
  RegisterFile RegisterFile_132 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_132_clock),
    .reset(RegisterFile_132_reset),
    .io_configuration(RegisterFile_132_io_configuration),
    .io_inputs_0(RegisterFile_132_io_inputs_0),
    .io_outs_0(RegisterFile_132_io_outs_0)
  );
  RegisterFile RegisterFile_133 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_133_clock),
    .reset(RegisterFile_133_reset),
    .io_configuration(RegisterFile_133_io_configuration),
    .io_inputs_0(RegisterFile_133_io_inputs_0),
    .io_outs_0(RegisterFile_133_io_outs_0)
  );
  RegisterFile RegisterFile_134 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_134_clock),
    .reset(RegisterFile_134_reset),
    .io_configuration(RegisterFile_134_io_configuration),
    .io_inputs_0(RegisterFile_134_io_inputs_0),
    .io_outs_0(RegisterFile_134_io_outs_0)
  );
  RegisterFile RegisterFile_135 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_135_clock),
    .reset(RegisterFile_135_reset),
    .io_configuration(RegisterFile_135_io_configuration),
    .io_inputs_0(RegisterFile_135_io_inputs_0),
    .io_outs_0(RegisterFile_135_io_outs_0)
  );
  RegisterFile RegisterFile_136 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_136_clock),
    .reset(RegisterFile_136_reset),
    .io_configuration(RegisterFile_136_io_configuration),
    .io_inputs_0(RegisterFile_136_io_inputs_0),
    .io_outs_0(RegisterFile_136_io_outs_0)
  );
  RegisterFile RegisterFile_137 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_137_clock),
    .reset(RegisterFile_137_reset),
    .io_configuration(RegisterFile_137_io_configuration),
    .io_inputs_0(RegisterFile_137_io_inputs_0),
    .io_outs_0(RegisterFile_137_io_outs_0)
  );
  RegisterFile RegisterFile_138 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_138_clock),
    .reset(RegisterFile_138_reset),
    .io_configuration(RegisterFile_138_io_configuration),
    .io_inputs_0(RegisterFile_138_io_inputs_0),
    .io_outs_0(RegisterFile_138_io_outs_0)
  );
  RegisterFile RegisterFile_139 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_139_clock),
    .reset(RegisterFile_139_reset),
    .io_configuration(RegisterFile_139_io_configuration),
    .io_inputs_0(RegisterFile_139_io_inputs_0),
    .io_outs_0(RegisterFile_139_io_outs_0)
  );
  RegisterFile RegisterFile_140 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_140_clock),
    .reset(RegisterFile_140_reset),
    .io_configuration(RegisterFile_140_io_configuration),
    .io_inputs_0(RegisterFile_140_io_inputs_0),
    .io_outs_0(RegisterFile_140_io_outs_0)
  );
  RegisterFile RegisterFile_141 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_141_clock),
    .reset(RegisterFile_141_reset),
    .io_configuration(RegisterFile_141_io_configuration),
    .io_inputs_0(RegisterFile_141_io_inputs_0),
    .io_outs_0(RegisterFile_141_io_outs_0)
  );
  RegisterFile RegisterFile_142 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_142_clock),
    .reset(RegisterFile_142_reset),
    .io_configuration(RegisterFile_142_io_configuration),
    .io_inputs_0(RegisterFile_142_io_inputs_0),
    .io_outs_0(RegisterFile_142_io_outs_0)
  );
  RegisterFile RegisterFile_143 ( // @[TopModule.scala 158:21]
    .clock(RegisterFile_143_clock),
    .reset(RegisterFile_143_reset),
    .io_configuration(RegisterFile_143_io_configuration),
    .io_inputs_0(RegisterFile_143_io_inputs_0),
    .io_outs_0(RegisterFile_143_io_outs_0)
  );
  Multiplexer Multiplexer ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_io_configuration),
    .io_inputs_4(Multiplexer_io_inputs_4),
    .io_inputs_3(Multiplexer_io_inputs_3),
    .io_inputs_2(Multiplexer_io_inputs_2),
    .io_inputs_1(Multiplexer_io_inputs_1),
    .io_inputs_0(Multiplexer_io_inputs_0),
    .io_outs_0(Multiplexer_io_outs_0)
  );
  Multiplexer Multiplexer_1 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_1_io_configuration),
    .io_inputs_4(Multiplexer_1_io_inputs_4),
    .io_inputs_3(Multiplexer_1_io_inputs_3),
    .io_inputs_2(Multiplexer_1_io_inputs_2),
    .io_inputs_1(Multiplexer_1_io_inputs_1),
    .io_inputs_0(Multiplexer_1_io_inputs_0),
    .io_outs_0(Multiplexer_1_io_outs_0)
  );
  Multiplexer Multiplexer_2 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_2_io_configuration),
    .io_inputs_4(Multiplexer_2_io_inputs_4),
    .io_inputs_3(Multiplexer_2_io_inputs_3),
    .io_inputs_2(Multiplexer_2_io_inputs_2),
    .io_inputs_1(Multiplexer_2_io_inputs_1),
    .io_inputs_0(Multiplexer_2_io_inputs_0),
    .io_outs_0(Multiplexer_2_io_outs_0)
  );
  Multiplexer Multiplexer_3 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_3_io_configuration),
    .io_inputs_4(Multiplexer_3_io_inputs_4),
    .io_inputs_3(Multiplexer_3_io_inputs_3),
    .io_inputs_2(Multiplexer_3_io_inputs_2),
    .io_inputs_1(Multiplexer_3_io_inputs_1),
    .io_inputs_0(Multiplexer_3_io_inputs_0),
    .io_outs_0(Multiplexer_3_io_outs_0)
  );
  Multiplexer Multiplexer_4 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_4_io_configuration),
    .io_inputs_4(Multiplexer_4_io_inputs_4),
    .io_inputs_3(Multiplexer_4_io_inputs_3),
    .io_inputs_2(Multiplexer_4_io_inputs_2),
    .io_inputs_1(Multiplexer_4_io_inputs_1),
    .io_inputs_0(Multiplexer_4_io_inputs_0),
    .io_outs_0(Multiplexer_4_io_outs_0)
  );
  Multiplexer_5 Multiplexer_5 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_5_io_configuration),
    .io_inputs_1(Multiplexer_5_io_inputs_1),
    .io_inputs_0(Multiplexer_5_io_inputs_0),
    .io_outs_0(Multiplexer_5_io_outs_0)
  );
  Multiplexer_5 Multiplexer_6 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_6_io_configuration),
    .io_inputs_1(Multiplexer_6_io_inputs_1),
    .io_inputs_0(Multiplexer_6_io_inputs_0),
    .io_outs_0(Multiplexer_6_io_outs_0)
  );
  Multiplexer_5 Multiplexer_7 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_7_io_configuration),
    .io_inputs_1(Multiplexer_7_io_inputs_1),
    .io_inputs_0(Multiplexer_7_io_inputs_0),
    .io_outs_0(Multiplexer_7_io_outs_0)
  );
  Multiplexer_8 Multiplexer_8 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_8_io_configuration),
    .io_inputs_5(Multiplexer_8_io_inputs_5),
    .io_inputs_4(Multiplexer_8_io_inputs_4),
    .io_inputs_3(Multiplexer_8_io_inputs_3),
    .io_inputs_2(Multiplexer_8_io_inputs_2),
    .io_inputs_1(Multiplexer_8_io_inputs_1),
    .io_inputs_0(Multiplexer_8_io_inputs_0),
    .io_outs_0(Multiplexer_8_io_outs_0)
  );
  Multiplexer_8 Multiplexer_9 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_9_io_configuration),
    .io_inputs_5(Multiplexer_9_io_inputs_5),
    .io_inputs_4(Multiplexer_9_io_inputs_4),
    .io_inputs_3(Multiplexer_9_io_inputs_3),
    .io_inputs_2(Multiplexer_9_io_inputs_2),
    .io_inputs_1(Multiplexer_9_io_inputs_1),
    .io_inputs_0(Multiplexer_9_io_inputs_0),
    .io_outs_0(Multiplexer_9_io_outs_0)
  );
  Multiplexer_8 Multiplexer_10 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_10_io_configuration),
    .io_inputs_5(Multiplexer_10_io_inputs_5),
    .io_inputs_4(Multiplexer_10_io_inputs_4),
    .io_inputs_3(Multiplexer_10_io_inputs_3),
    .io_inputs_2(Multiplexer_10_io_inputs_2),
    .io_inputs_1(Multiplexer_10_io_inputs_1),
    .io_inputs_0(Multiplexer_10_io_inputs_0),
    .io_outs_0(Multiplexer_10_io_outs_0)
  );
  Multiplexer_8 Multiplexer_11 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_11_io_configuration),
    .io_inputs_5(Multiplexer_11_io_inputs_5),
    .io_inputs_4(Multiplexer_11_io_inputs_4),
    .io_inputs_3(Multiplexer_11_io_inputs_3),
    .io_inputs_2(Multiplexer_11_io_inputs_2),
    .io_inputs_1(Multiplexer_11_io_inputs_1),
    .io_inputs_0(Multiplexer_11_io_inputs_0),
    .io_outs_0(Multiplexer_11_io_outs_0)
  );
  Multiplexer_8 Multiplexer_12 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_12_io_configuration),
    .io_inputs_5(Multiplexer_12_io_inputs_5),
    .io_inputs_4(Multiplexer_12_io_inputs_4),
    .io_inputs_3(Multiplexer_12_io_inputs_3),
    .io_inputs_2(Multiplexer_12_io_inputs_2),
    .io_inputs_1(Multiplexer_12_io_inputs_1),
    .io_inputs_0(Multiplexer_12_io_inputs_0),
    .io_outs_0(Multiplexer_12_io_outs_0)
  );
  Multiplexer_8 Multiplexer_13 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_13_io_configuration),
    .io_inputs_5(Multiplexer_13_io_inputs_5),
    .io_inputs_4(Multiplexer_13_io_inputs_4),
    .io_inputs_3(Multiplexer_13_io_inputs_3),
    .io_inputs_2(Multiplexer_13_io_inputs_2),
    .io_inputs_1(Multiplexer_13_io_inputs_1),
    .io_inputs_0(Multiplexer_13_io_inputs_0),
    .io_outs_0(Multiplexer_13_io_outs_0)
  );
  Multiplexer_5 Multiplexer_14 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_14_io_configuration),
    .io_inputs_1(Multiplexer_14_io_inputs_1),
    .io_inputs_0(Multiplexer_14_io_inputs_0),
    .io_outs_0(Multiplexer_14_io_outs_0)
  );
  Multiplexer_5 Multiplexer_15 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_15_io_configuration),
    .io_inputs_1(Multiplexer_15_io_inputs_1),
    .io_inputs_0(Multiplexer_15_io_inputs_0),
    .io_outs_0(Multiplexer_15_io_outs_0)
  );
  Multiplexer_5 Multiplexer_16 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_16_io_configuration),
    .io_inputs_1(Multiplexer_16_io_inputs_1),
    .io_inputs_0(Multiplexer_16_io_inputs_0),
    .io_outs_0(Multiplexer_16_io_outs_0)
  );
  Multiplexer_5 Multiplexer_17 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_17_io_configuration),
    .io_inputs_1(Multiplexer_17_io_inputs_1),
    .io_inputs_0(Multiplexer_17_io_inputs_0),
    .io_outs_0(Multiplexer_17_io_outs_0)
  );
  Multiplexer_8 Multiplexer_18 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_18_io_configuration),
    .io_inputs_5(Multiplexer_18_io_inputs_5),
    .io_inputs_4(Multiplexer_18_io_inputs_4),
    .io_inputs_3(Multiplexer_18_io_inputs_3),
    .io_inputs_2(Multiplexer_18_io_inputs_2),
    .io_inputs_1(Multiplexer_18_io_inputs_1),
    .io_inputs_0(Multiplexer_18_io_inputs_0),
    .io_outs_0(Multiplexer_18_io_outs_0)
  );
  Multiplexer_8 Multiplexer_19 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_19_io_configuration),
    .io_inputs_5(Multiplexer_19_io_inputs_5),
    .io_inputs_4(Multiplexer_19_io_inputs_4),
    .io_inputs_3(Multiplexer_19_io_inputs_3),
    .io_inputs_2(Multiplexer_19_io_inputs_2),
    .io_inputs_1(Multiplexer_19_io_inputs_1),
    .io_inputs_0(Multiplexer_19_io_inputs_0),
    .io_outs_0(Multiplexer_19_io_outs_0)
  );
  Multiplexer_8 Multiplexer_20 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_20_io_configuration),
    .io_inputs_5(Multiplexer_20_io_inputs_5),
    .io_inputs_4(Multiplexer_20_io_inputs_4),
    .io_inputs_3(Multiplexer_20_io_inputs_3),
    .io_inputs_2(Multiplexer_20_io_inputs_2),
    .io_inputs_1(Multiplexer_20_io_inputs_1),
    .io_inputs_0(Multiplexer_20_io_inputs_0),
    .io_outs_0(Multiplexer_20_io_outs_0)
  );
  Multiplexer_8 Multiplexer_21 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_21_io_configuration),
    .io_inputs_5(Multiplexer_21_io_inputs_5),
    .io_inputs_4(Multiplexer_21_io_inputs_4),
    .io_inputs_3(Multiplexer_21_io_inputs_3),
    .io_inputs_2(Multiplexer_21_io_inputs_2),
    .io_inputs_1(Multiplexer_21_io_inputs_1),
    .io_inputs_0(Multiplexer_21_io_inputs_0),
    .io_outs_0(Multiplexer_21_io_outs_0)
  );
  Multiplexer_8 Multiplexer_22 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_22_io_configuration),
    .io_inputs_5(Multiplexer_22_io_inputs_5),
    .io_inputs_4(Multiplexer_22_io_inputs_4),
    .io_inputs_3(Multiplexer_22_io_inputs_3),
    .io_inputs_2(Multiplexer_22_io_inputs_2),
    .io_inputs_1(Multiplexer_22_io_inputs_1),
    .io_inputs_0(Multiplexer_22_io_inputs_0),
    .io_outs_0(Multiplexer_22_io_outs_0)
  );
  Multiplexer_8 Multiplexer_23 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_23_io_configuration),
    .io_inputs_5(Multiplexer_23_io_inputs_5),
    .io_inputs_4(Multiplexer_23_io_inputs_4),
    .io_inputs_3(Multiplexer_23_io_inputs_3),
    .io_inputs_2(Multiplexer_23_io_inputs_2),
    .io_inputs_1(Multiplexer_23_io_inputs_1),
    .io_inputs_0(Multiplexer_23_io_inputs_0),
    .io_outs_0(Multiplexer_23_io_outs_0)
  );
  Multiplexer_5 Multiplexer_24 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_24_io_configuration),
    .io_inputs_1(Multiplexer_24_io_inputs_1),
    .io_inputs_0(Multiplexer_24_io_inputs_0),
    .io_outs_0(Multiplexer_24_io_outs_0)
  );
  Multiplexer_5 Multiplexer_25 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_25_io_configuration),
    .io_inputs_1(Multiplexer_25_io_inputs_1),
    .io_inputs_0(Multiplexer_25_io_inputs_0),
    .io_outs_0(Multiplexer_25_io_outs_0)
  );
  Multiplexer_5 Multiplexer_26 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_26_io_configuration),
    .io_inputs_1(Multiplexer_26_io_inputs_1),
    .io_inputs_0(Multiplexer_26_io_inputs_0),
    .io_outs_0(Multiplexer_26_io_outs_0)
  );
  Multiplexer_5 Multiplexer_27 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_27_io_configuration),
    .io_inputs_1(Multiplexer_27_io_inputs_1),
    .io_inputs_0(Multiplexer_27_io_inputs_0),
    .io_outs_0(Multiplexer_27_io_outs_0)
  );
  Multiplexer_8 Multiplexer_28 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_28_io_configuration),
    .io_inputs_5(Multiplexer_28_io_inputs_5),
    .io_inputs_4(Multiplexer_28_io_inputs_4),
    .io_inputs_3(Multiplexer_28_io_inputs_3),
    .io_inputs_2(Multiplexer_28_io_inputs_2),
    .io_inputs_1(Multiplexer_28_io_inputs_1),
    .io_inputs_0(Multiplexer_28_io_inputs_0),
    .io_outs_0(Multiplexer_28_io_outs_0)
  );
  Multiplexer_8 Multiplexer_29 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_29_io_configuration),
    .io_inputs_5(Multiplexer_29_io_inputs_5),
    .io_inputs_4(Multiplexer_29_io_inputs_4),
    .io_inputs_3(Multiplexer_29_io_inputs_3),
    .io_inputs_2(Multiplexer_29_io_inputs_2),
    .io_inputs_1(Multiplexer_29_io_inputs_1),
    .io_inputs_0(Multiplexer_29_io_inputs_0),
    .io_outs_0(Multiplexer_29_io_outs_0)
  );
  Multiplexer_8 Multiplexer_30 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_30_io_configuration),
    .io_inputs_5(Multiplexer_30_io_inputs_5),
    .io_inputs_4(Multiplexer_30_io_inputs_4),
    .io_inputs_3(Multiplexer_30_io_inputs_3),
    .io_inputs_2(Multiplexer_30_io_inputs_2),
    .io_inputs_1(Multiplexer_30_io_inputs_1),
    .io_inputs_0(Multiplexer_30_io_inputs_0),
    .io_outs_0(Multiplexer_30_io_outs_0)
  );
  Multiplexer_8 Multiplexer_31 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_31_io_configuration),
    .io_inputs_5(Multiplexer_31_io_inputs_5),
    .io_inputs_4(Multiplexer_31_io_inputs_4),
    .io_inputs_3(Multiplexer_31_io_inputs_3),
    .io_inputs_2(Multiplexer_31_io_inputs_2),
    .io_inputs_1(Multiplexer_31_io_inputs_1),
    .io_inputs_0(Multiplexer_31_io_inputs_0),
    .io_outs_0(Multiplexer_31_io_outs_0)
  );
  Multiplexer_8 Multiplexer_32 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_32_io_configuration),
    .io_inputs_5(Multiplexer_32_io_inputs_5),
    .io_inputs_4(Multiplexer_32_io_inputs_4),
    .io_inputs_3(Multiplexer_32_io_inputs_3),
    .io_inputs_2(Multiplexer_32_io_inputs_2),
    .io_inputs_1(Multiplexer_32_io_inputs_1),
    .io_inputs_0(Multiplexer_32_io_inputs_0),
    .io_outs_0(Multiplexer_32_io_outs_0)
  );
  Multiplexer_8 Multiplexer_33 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_33_io_configuration),
    .io_inputs_5(Multiplexer_33_io_inputs_5),
    .io_inputs_4(Multiplexer_33_io_inputs_4),
    .io_inputs_3(Multiplexer_33_io_inputs_3),
    .io_inputs_2(Multiplexer_33_io_inputs_2),
    .io_inputs_1(Multiplexer_33_io_inputs_1),
    .io_inputs_0(Multiplexer_33_io_inputs_0),
    .io_outs_0(Multiplexer_33_io_outs_0)
  );
  Multiplexer_5 Multiplexer_34 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_34_io_configuration),
    .io_inputs_1(Multiplexer_34_io_inputs_1),
    .io_inputs_0(Multiplexer_34_io_inputs_0),
    .io_outs_0(Multiplexer_34_io_outs_0)
  );
  Multiplexer_5 Multiplexer_35 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_35_io_configuration),
    .io_inputs_1(Multiplexer_35_io_inputs_1),
    .io_inputs_0(Multiplexer_35_io_inputs_0),
    .io_outs_0(Multiplexer_35_io_outs_0)
  );
  Multiplexer_5 Multiplexer_36 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_36_io_configuration),
    .io_inputs_1(Multiplexer_36_io_inputs_1),
    .io_inputs_0(Multiplexer_36_io_inputs_0),
    .io_outs_0(Multiplexer_36_io_outs_0)
  );
  Multiplexer_5 Multiplexer_37 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_37_io_configuration),
    .io_inputs_1(Multiplexer_37_io_inputs_1),
    .io_inputs_0(Multiplexer_37_io_inputs_0),
    .io_outs_0(Multiplexer_37_io_outs_0)
  );
  Multiplexer_8 Multiplexer_38 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_38_io_configuration),
    .io_inputs_5(Multiplexer_38_io_inputs_5),
    .io_inputs_4(Multiplexer_38_io_inputs_4),
    .io_inputs_3(Multiplexer_38_io_inputs_3),
    .io_inputs_2(Multiplexer_38_io_inputs_2),
    .io_inputs_1(Multiplexer_38_io_inputs_1),
    .io_inputs_0(Multiplexer_38_io_inputs_0),
    .io_outs_0(Multiplexer_38_io_outs_0)
  );
  Multiplexer_8 Multiplexer_39 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_39_io_configuration),
    .io_inputs_5(Multiplexer_39_io_inputs_5),
    .io_inputs_4(Multiplexer_39_io_inputs_4),
    .io_inputs_3(Multiplexer_39_io_inputs_3),
    .io_inputs_2(Multiplexer_39_io_inputs_2),
    .io_inputs_1(Multiplexer_39_io_inputs_1),
    .io_inputs_0(Multiplexer_39_io_inputs_0),
    .io_outs_0(Multiplexer_39_io_outs_0)
  );
  Multiplexer_8 Multiplexer_40 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_40_io_configuration),
    .io_inputs_5(Multiplexer_40_io_inputs_5),
    .io_inputs_4(Multiplexer_40_io_inputs_4),
    .io_inputs_3(Multiplexer_40_io_inputs_3),
    .io_inputs_2(Multiplexer_40_io_inputs_2),
    .io_inputs_1(Multiplexer_40_io_inputs_1),
    .io_inputs_0(Multiplexer_40_io_inputs_0),
    .io_outs_0(Multiplexer_40_io_outs_0)
  );
  Multiplexer_8 Multiplexer_41 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_41_io_configuration),
    .io_inputs_5(Multiplexer_41_io_inputs_5),
    .io_inputs_4(Multiplexer_41_io_inputs_4),
    .io_inputs_3(Multiplexer_41_io_inputs_3),
    .io_inputs_2(Multiplexer_41_io_inputs_2),
    .io_inputs_1(Multiplexer_41_io_inputs_1),
    .io_inputs_0(Multiplexer_41_io_inputs_0),
    .io_outs_0(Multiplexer_41_io_outs_0)
  );
  Multiplexer_8 Multiplexer_42 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_42_io_configuration),
    .io_inputs_5(Multiplexer_42_io_inputs_5),
    .io_inputs_4(Multiplexer_42_io_inputs_4),
    .io_inputs_3(Multiplexer_42_io_inputs_3),
    .io_inputs_2(Multiplexer_42_io_inputs_2),
    .io_inputs_1(Multiplexer_42_io_inputs_1),
    .io_inputs_0(Multiplexer_42_io_inputs_0),
    .io_outs_0(Multiplexer_42_io_outs_0)
  );
  Multiplexer_8 Multiplexer_43 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_43_io_configuration),
    .io_inputs_5(Multiplexer_43_io_inputs_5),
    .io_inputs_4(Multiplexer_43_io_inputs_4),
    .io_inputs_3(Multiplexer_43_io_inputs_3),
    .io_inputs_2(Multiplexer_43_io_inputs_2),
    .io_inputs_1(Multiplexer_43_io_inputs_1),
    .io_inputs_0(Multiplexer_43_io_inputs_0),
    .io_outs_0(Multiplexer_43_io_outs_0)
  );
  Multiplexer_5 Multiplexer_44 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_44_io_configuration),
    .io_inputs_1(Multiplexer_44_io_inputs_1),
    .io_inputs_0(Multiplexer_44_io_inputs_0),
    .io_outs_0(Multiplexer_44_io_outs_0)
  );
  Multiplexer_5 Multiplexer_45 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_45_io_configuration),
    .io_inputs_1(Multiplexer_45_io_inputs_1),
    .io_inputs_0(Multiplexer_45_io_inputs_0),
    .io_outs_0(Multiplexer_45_io_outs_0)
  );
  Multiplexer_5 Multiplexer_46 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_46_io_configuration),
    .io_inputs_1(Multiplexer_46_io_inputs_1),
    .io_inputs_0(Multiplexer_46_io_inputs_0),
    .io_outs_0(Multiplexer_46_io_outs_0)
  );
  Multiplexer_5 Multiplexer_47 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_47_io_configuration),
    .io_inputs_1(Multiplexer_47_io_inputs_1),
    .io_inputs_0(Multiplexer_47_io_inputs_0),
    .io_outs_0(Multiplexer_47_io_outs_0)
  );
  Multiplexer Multiplexer_48 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_48_io_configuration),
    .io_inputs_4(Multiplexer_48_io_inputs_4),
    .io_inputs_3(Multiplexer_48_io_inputs_3),
    .io_inputs_2(Multiplexer_48_io_inputs_2),
    .io_inputs_1(Multiplexer_48_io_inputs_1),
    .io_inputs_0(Multiplexer_48_io_inputs_0),
    .io_outs_0(Multiplexer_48_io_outs_0)
  );
  Multiplexer Multiplexer_49 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_49_io_configuration),
    .io_inputs_4(Multiplexer_49_io_inputs_4),
    .io_inputs_3(Multiplexer_49_io_inputs_3),
    .io_inputs_2(Multiplexer_49_io_inputs_2),
    .io_inputs_1(Multiplexer_49_io_inputs_1),
    .io_inputs_0(Multiplexer_49_io_inputs_0),
    .io_outs_0(Multiplexer_49_io_outs_0)
  );
  Multiplexer Multiplexer_50 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_50_io_configuration),
    .io_inputs_4(Multiplexer_50_io_inputs_4),
    .io_inputs_3(Multiplexer_50_io_inputs_3),
    .io_inputs_2(Multiplexer_50_io_inputs_2),
    .io_inputs_1(Multiplexer_50_io_inputs_1),
    .io_inputs_0(Multiplexer_50_io_inputs_0),
    .io_outs_0(Multiplexer_50_io_outs_0)
  );
  Multiplexer Multiplexer_51 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_51_io_configuration),
    .io_inputs_4(Multiplexer_51_io_inputs_4),
    .io_inputs_3(Multiplexer_51_io_inputs_3),
    .io_inputs_2(Multiplexer_51_io_inputs_2),
    .io_inputs_1(Multiplexer_51_io_inputs_1),
    .io_inputs_0(Multiplexer_51_io_inputs_0),
    .io_outs_0(Multiplexer_51_io_outs_0)
  );
  Multiplexer Multiplexer_52 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_52_io_configuration),
    .io_inputs_4(Multiplexer_52_io_inputs_4),
    .io_inputs_3(Multiplexer_52_io_inputs_3),
    .io_inputs_2(Multiplexer_52_io_inputs_2),
    .io_inputs_1(Multiplexer_52_io_inputs_1),
    .io_inputs_0(Multiplexer_52_io_inputs_0),
    .io_outs_0(Multiplexer_52_io_outs_0)
  );
  Multiplexer_5 Multiplexer_53 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_53_io_configuration),
    .io_inputs_1(Multiplexer_53_io_inputs_1),
    .io_inputs_0(Multiplexer_53_io_inputs_0),
    .io_outs_0(Multiplexer_53_io_outs_0)
  );
  Multiplexer_5 Multiplexer_54 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_54_io_configuration),
    .io_inputs_1(Multiplexer_54_io_inputs_1),
    .io_inputs_0(Multiplexer_54_io_inputs_0),
    .io_outs_0(Multiplexer_54_io_outs_0)
  );
  Multiplexer_5 Multiplexer_55 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_55_io_configuration),
    .io_inputs_1(Multiplexer_55_io_inputs_1),
    .io_inputs_0(Multiplexer_55_io_inputs_0),
    .io_outs_0(Multiplexer_55_io_outs_0)
  );
  Multiplexer Multiplexer_56 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_56_io_configuration),
    .io_inputs_4(Multiplexer_56_io_inputs_4),
    .io_inputs_3(Multiplexer_56_io_inputs_3),
    .io_inputs_2(Multiplexer_56_io_inputs_2),
    .io_inputs_1(Multiplexer_56_io_inputs_1),
    .io_inputs_0(Multiplexer_56_io_inputs_0),
    .io_outs_0(Multiplexer_56_io_outs_0)
  );
  Multiplexer Multiplexer_57 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_57_io_configuration),
    .io_inputs_4(Multiplexer_57_io_inputs_4),
    .io_inputs_3(Multiplexer_57_io_inputs_3),
    .io_inputs_2(Multiplexer_57_io_inputs_2),
    .io_inputs_1(Multiplexer_57_io_inputs_1),
    .io_inputs_0(Multiplexer_57_io_inputs_0),
    .io_outs_0(Multiplexer_57_io_outs_0)
  );
  Multiplexer Multiplexer_58 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_58_io_configuration),
    .io_inputs_4(Multiplexer_58_io_inputs_4),
    .io_inputs_3(Multiplexer_58_io_inputs_3),
    .io_inputs_2(Multiplexer_58_io_inputs_2),
    .io_inputs_1(Multiplexer_58_io_inputs_1),
    .io_inputs_0(Multiplexer_58_io_inputs_0),
    .io_outs_0(Multiplexer_58_io_outs_0)
  );
  Multiplexer Multiplexer_59 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_59_io_configuration),
    .io_inputs_4(Multiplexer_59_io_inputs_4),
    .io_inputs_3(Multiplexer_59_io_inputs_3),
    .io_inputs_2(Multiplexer_59_io_inputs_2),
    .io_inputs_1(Multiplexer_59_io_inputs_1),
    .io_inputs_0(Multiplexer_59_io_inputs_0),
    .io_outs_0(Multiplexer_59_io_outs_0)
  );
  Multiplexer Multiplexer_60 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_60_io_configuration),
    .io_inputs_4(Multiplexer_60_io_inputs_4),
    .io_inputs_3(Multiplexer_60_io_inputs_3),
    .io_inputs_2(Multiplexer_60_io_inputs_2),
    .io_inputs_1(Multiplexer_60_io_inputs_1),
    .io_inputs_0(Multiplexer_60_io_inputs_0),
    .io_outs_0(Multiplexer_60_io_outs_0)
  );
  Multiplexer_5 Multiplexer_61 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_61_io_configuration),
    .io_inputs_1(Multiplexer_61_io_inputs_1),
    .io_inputs_0(Multiplexer_61_io_inputs_0),
    .io_outs_0(Multiplexer_61_io_outs_0)
  );
  Multiplexer_5 Multiplexer_62 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_62_io_configuration),
    .io_inputs_1(Multiplexer_62_io_inputs_1),
    .io_inputs_0(Multiplexer_62_io_inputs_0),
    .io_outs_0(Multiplexer_62_io_outs_0)
  );
  Multiplexer_5 Multiplexer_63 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_63_io_configuration),
    .io_inputs_1(Multiplexer_63_io_inputs_1),
    .io_inputs_0(Multiplexer_63_io_inputs_0),
    .io_outs_0(Multiplexer_63_io_outs_0)
  );
  Multiplexer_8 Multiplexer_64 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_64_io_configuration),
    .io_inputs_5(Multiplexer_64_io_inputs_5),
    .io_inputs_4(Multiplexer_64_io_inputs_4),
    .io_inputs_3(Multiplexer_64_io_inputs_3),
    .io_inputs_2(Multiplexer_64_io_inputs_2),
    .io_inputs_1(Multiplexer_64_io_inputs_1),
    .io_inputs_0(Multiplexer_64_io_inputs_0),
    .io_outs_0(Multiplexer_64_io_outs_0)
  );
  Multiplexer_8 Multiplexer_65 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_65_io_configuration),
    .io_inputs_5(Multiplexer_65_io_inputs_5),
    .io_inputs_4(Multiplexer_65_io_inputs_4),
    .io_inputs_3(Multiplexer_65_io_inputs_3),
    .io_inputs_2(Multiplexer_65_io_inputs_2),
    .io_inputs_1(Multiplexer_65_io_inputs_1),
    .io_inputs_0(Multiplexer_65_io_inputs_0),
    .io_outs_0(Multiplexer_65_io_outs_0)
  );
  Multiplexer_8 Multiplexer_66 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_66_io_configuration),
    .io_inputs_5(Multiplexer_66_io_inputs_5),
    .io_inputs_4(Multiplexer_66_io_inputs_4),
    .io_inputs_3(Multiplexer_66_io_inputs_3),
    .io_inputs_2(Multiplexer_66_io_inputs_2),
    .io_inputs_1(Multiplexer_66_io_inputs_1),
    .io_inputs_0(Multiplexer_66_io_inputs_0),
    .io_outs_0(Multiplexer_66_io_outs_0)
  );
  Multiplexer_8 Multiplexer_67 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_67_io_configuration),
    .io_inputs_5(Multiplexer_67_io_inputs_5),
    .io_inputs_4(Multiplexer_67_io_inputs_4),
    .io_inputs_3(Multiplexer_67_io_inputs_3),
    .io_inputs_2(Multiplexer_67_io_inputs_2),
    .io_inputs_1(Multiplexer_67_io_inputs_1),
    .io_inputs_0(Multiplexer_67_io_inputs_0),
    .io_outs_0(Multiplexer_67_io_outs_0)
  );
  Multiplexer_8 Multiplexer_68 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_68_io_configuration),
    .io_inputs_5(Multiplexer_68_io_inputs_5),
    .io_inputs_4(Multiplexer_68_io_inputs_4),
    .io_inputs_3(Multiplexer_68_io_inputs_3),
    .io_inputs_2(Multiplexer_68_io_inputs_2),
    .io_inputs_1(Multiplexer_68_io_inputs_1),
    .io_inputs_0(Multiplexer_68_io_inputs_0),
    .io_outs_0(Multiplexer_68_io_outs_0)
  );
  Multiplexer_8 Multiplexer_69 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_69_io_configuration),
    .io_inputs_5(Multiplexer_69_io_inputs_5),
    .io_inputs_4(Multiplexer_69_io_inputs_4),
    .io_inputs_3(Multiplexer_69_io_inputs_3),
    .io_inputs_2(Multiplexer_69_io_inputs_2),
    .io_inputs_1(Multiplexer_69_io_inputs_1),
    .io_inputs_0(Multiplexer_69_io_inputs_0),
    .io_outs_0(Multiplexer_69_io_outs_0)
  );
  Multiplexer_5 Multiplexer_70 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_70_io_configuration),
    .io_inputs_1(Multiplexer_70_io_inputs_1),
    .io_inputs_0(Multiplexer_70_io_inputs_0),
    .io_outs_0(Multiplexer_70_io_outs_0)
  );
  Multiplexer_5 Multiplexer_71 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_71_io_configuration),
    .io_inputs_1(Multiplexer_71_io_inputs_1),
    .io_inputs_0(Multiplexer_71_io_inputs_0),
    .io_outs_0(Multiplexer_71_io_outs_0)
  );
  Multiplexer_5 Multiplexer_72 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_72_io_configuration),
    .io_inputs_1(Multiplexer_72_io_inputs_1),
    .io_inputs_0(Multiplexer_72_io_inputs_0),
    .io_outs_0(Multiplexer_72_io_outs_0)
  );
  Multiplexer_5 Multiplexer_73 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_73_io_configuration),
    .io_inputs_1(Multiplexer_73_io_inputs_1),
    .io_inputs_0(Multiplexer_73_io_inputs_0),
    .io_outs_0(Multiplexer_73_io_outs_0)
  );
  Multiplexer_8 Multiplexer_74 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_74_io_configuration),
    .io_inputs_5(Multiplexer_74_io_inputs_5),
    .io_inputs_4(Multiplexer_74_io_inputs_4),
    .io_inputs_3(Multiplexer_74_io_inputs_3),
    .io_inputs_2(Multiplexer_74_io_inputs_2),
    .io_inputs_1(Multiplexer_74_io_inputs_1),
    .io_inputs_0(Multiplexer_74_io_inputs_0),
    .io_outs_0(Multiplexer_74_io_outs_0)
  );
  Multiplexer_8 Multiplexer_75 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_75_io_configuration),
    .io_inputs_5(Multiplexer_75_io_inputs_5),
    .io_inputs_4(Multiplexer_75_io_inputs_4),
    .io_inputs_3(Multiplexer_75_io_inputs_3),
    .io_inputs_2(Multiplexer_75_io_inputs_2),
    .io_inputs_1(Multiplexer_75_io_inputs_1),
    .io_inputs_0(Multiplexer_75_io_inputs_0),
    .io_outs_0(Multiplexer_75_io_outs_0)
  );
  Multiplexer_8 Multiplexer_76 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_76_io_configuration),
    .io_inputs_5(Multiplexer_76_io_inputs_5),
    .io_inputs_4(Multiplexer_76_io_inputs_4),
    .io_inputs_3(Multiplexer_76_io_inputs_3),
    .io_inputs_2(Multiplexer_76_io_inputs_2),
    .io_inputs_1(Multiplexer_76_io_inputs_1),
    .io_inputs_0(Multiplexer_76_io_inputs_0),
    .io_outs_0(Multiplexer_76_io_outs_0)
  );
  Multiplexer_8 Multiplexer_77 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_77_io_configuration),
    .io_inputs_5(Multiplexer_77_io_inputs_5),
    .io_inputs_4(Multiplexer_77_io_inputs_4),
    .io_inputs_3(Multiplexer_77_io_inputs_3),
    .io_inputs_2(Multiplexer_77_io_inputs_2),
    .io_inputs_1(Multiplexer_77_io_inputs_1),
    .io_inputs_0(Multiplexer_77_io_inputs_0),
    .io_outs_0(Multiplexer_77_io_outs_0)
  );
  Multiplexer_8 Multiplexer_78 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_78_io_configuration),
    .io_inputs_5(Multiplexer_78_io_inputs_5),
    .io_inputs_4(Multiplexer_78_io_inputs_4),
    .io_inputs_3(Multiplexer_78_io_inputs_3),
    .io_inputs_2(Multiplexer_78_io_inputs_2),
    .io_inputs_1(Multiplexer_78_io_inputs_1),
    .io_inputs_0(Multiplexer_78_io_inputs_0),
    .io_outs_0(Multiplexer_78_io_outs_0)
  );
  Multiplexer_8 Multiplexer_79 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_79_io_configuration),
    .io_inputs_5(Multiplexer_79_io_inputs_5),
    .io_inputs_4(Multiplexer_79_io_inputs_4),
    .io_inputs_3(Multiplexer_79_io_inputs_3),
    .io_inputs_2(Multiplexer_79_io_inputs_2),
    .io_inputs_1(Multiplexer_79_io_inputs_1),
    .io_inputs_0(Multiplexer_79_io_inputs_0),
    .io_outs_0(Multiplexer_79_io_outs_0)
  );
  Multiplexer_5 Multiplexer_80 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_80_io_configuration),
    .io_inputs_1(Multiplexer_80_io_inputs_1),
    .io_inputs_0(Multiplexer_80_io_inputs_0),
    .io_outs_0(Multiplexer_80_io_outs_0)
  );
  Multiplexer_5 Multiplexer_81 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_81_io_configuration),
    .io_inputs_1(Multiplexer_81_io_inputs_1),
    .io_inputs_0(Multiplexer_81_io_inputs_0),
    .io_outs_0(Multiplexer_81_io_outs_0)
  );
  Multiplexer_5 Multiplexer_82 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_82_io_configuration),
    .io_inputs_1(Multiplexer_82_io_inputs_1),
    .io_inputs_0(Multiplexer_82_io_inputs_0),
    .io_outs_0(Multiplexer_82_io_outs_0)
  );
  Multiplexer_5 Multiplexer_83 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_83_io_configuration),
    .io_inputs_1(Multiplexer_83_io_inputs_1),
    .io_inputs_0(Multiplexer_83_io_inputs_0),
    .io_outs_0(Multiplexer_83_io_outs_0)
  );
  Multiplexer_8 Multiplexer_84 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_84_io_configuration),
    .io_inputs_5(Multiplexer_84_io_inputs_5),
    .io_inputs_4(Multiplexer_84_io_inputs_4),
    .io_inputs_3(Multiplexer_84_io_inputs_3),
    .io_inputs_2(Multiplexer_84_io_inputs_2),
    .io_inputs_1(Multiplexer_84_io_inputs_1),
    .io_inputs_0(Multiplexer_84_io_inputs_0),
    .io_outs_0(Multiplexer_84_io_outs_0)
  );
  Multiplexer_8 Multiplexer_85 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_85_io_configuration),
    .io_inputs_5(Multiplexer_85_io_inputs_5),
    .io_inputs_4(Multiplexer_85_io_inputs_4),
    .io_inputs_3(Multiplexer_85_io_inputs_3),
    .io_inputs_2(Multiplexer_85_io_inputs_2),
    .io_inputs_1(Multiplexer_85_io_inputs_1),
    .io_inputs_0(Multiplexer_85_io_inputs_0),
    .io_outs_0(Multiplexer_85_io_outs_0)
  );
  Multiplexer_8 Multiplexer_86 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_86_io_configuration),
    .io_inputs_5(Multiplexer_86_io_inputs_5),
    .io_inputs_4(Multiplexer_86_io_inputs_4),
    .io_inputs_3(Multiplexer_86_io_inputs_3),
    .io_inputs_2(Multiplexer_86_io_inputs_2),
    .io_inputs_1(Multiplexer_86_io_inputs_1),
    .io_inputs_0(Multiplexer_86_io_inputs_0),
    .io_outs_0(Multiplexer_86_io_outs_0)
  );
  Multiplexer_8 Multiplexer_87 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_87_io_configuration),
    .io_inputs_5(Multiplexer_87_io_inputs_5),
    .io_inputs_4(Multiplexer_87_io_inputs_4),
    .io_inputs_3(Multiplexer_87_io_inputs_3),
    .io_inputs_2(Multiplexer_87_io_inputs_2),
    .io_inputs_1(Multiplexer_87_io_inputs_1),
    .io_inputs_0(Multiplexer_87_io_inputs_0),
    .io_outs_0(Multiplexer_87_io_outs_0)
  );
  Multiplexer_8 Multiplexer_88 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_88_io_configuration),
    .io_inputs_5(Multiplexer_88_io_inputs_5),
    .io_inputs_4(Multiplexer_88_io_inputs_4),
    .io_inputs_3(Multiplexer_88_io_inputs_3),
    .io_inputs_2(Multiplexer_88_io_inputs_2),
    .io_inputs_1(Multiplexer_88_io_inputs_1),
    .io_inputs_0(Multiplexer_88_io_inputs_0),
    .io_outs_0(Multiplexer_88_io_outs_0)
  );
  Multiplexer_8 Multiplexer_89 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_89_io_configuration),
    .io_inputs_5(Multiplexer_89_io_inputs_5),
    .io_inputs_4(Multiplexer_89_io_inputs_4),
    .io_inputs_3(Multiplexer_89_io_inputs_3),
    .io_inputs_2(Multiplexer_89_io_inputs_2),
    .io_inputs_1(Multiplexer_89_io_inputs_1),
    .io_inputs_0(Multiplexer_89_io_inputs_0),
    .io_outs_0(Multiplexer_89_io_outs_0)
  );
  Multiplexer_5 Multiplexer_90 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_90_io_configuration),
    .io_inputs_1(Multiplexer_90_io_inputs_1),
    .io_inputs_0(Multiplexer_90_io_inputs_0),
    .io_outs_0(Multiplexer_90_io_outs_0)
  );
  Multiplexer_5 Multiplexer_91 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_91_io_configuration),
    .io_inputs_1(Multiplexer_91_io_inputs_1),
    .io_inputs_0(Multiplexer_91_io_inputs_0),
    .io_outs_0(Multiplexer_91_io_outs_0)
  );
  Multiplexer_5 Multiplexer_92 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_92_io_configuration),
    .io_inputs_1(Multiplexer_92_io_inputs_1),
    .io_inputs_0(Multiplexer_92_io_inputs_0),
    .io_outs_0(Multiplexer_92_io_outs_0)
  );
  Multiplexer_5 Multiplexer_93 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_93_io_configuration),
    .io_inputs_1(Multiplexer_93_io_inputs_1),
    .io_inputs_0(Multiplexer_93_io_inputs_0),
    .io_outs_0(Multiplexer_93_io_outs_0)
  );
  Multiplexer_8 Multiplexer_94 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_94_io_configuration),
    .io_inputs_5(Multiplexer_94_io_inputs_5),
    .io_inputs_4(Multiplexer_94_io_inputs_4),
    .io_inputs_3(Multiplexer_94_io_inputs_3),
    .io_inputs_2(Multiplexer_94_io_inputs_2),
    .io_inputs_1(Multiplexer_94_io_inputs_1),
    .io_inputs_0(Multiplexer_94_io_inputs_0),
    .io_outs_0(Multiplexer_94_io_outs_0)
  );
  Multiplexer_8 Multiplexer_95 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_95_io_configuration),
    .io_inputs_5(Multiplexer_95_io_inputs_5),
    .io_inputs_4(Multiplexer_95_io_inputs_4),
    .io_inputs_3(Multiplexer_95_io_inputs_3),
    .io_inputs_2(Multiplexer_95_io_inputs_2),
    .io_inputs_1(Multiplexer_95_io_inputs_1),
    .io_inputs_0(Multiplexer_95_io_inputs_0),
    .io_outs_0(Multiplexer_95_io_outs_0)
  );
  Multiplexer_8 Multiplexer_96 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_96_io_configuration),
    .io_inputs_5(Multiplexer_96_io_inputs_5),
    .io_inputs_4(Multiplexer_96_io_inputs_4),
    .io_inputs_3(Multiplexer_96_io_inputs_3),
    .io_inputs_2(Multiplexer_96_io_inputs_2),
    .io_inputs_1(Multiplexer_96_io_inputs_1),
    .io_inputs_0(Multiplexer_96_io_inputs_0),
    .io_outs_0(Multiplexer_96_io_outs_0)
  );
  Multiplexer_8 Multiplexer_97 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_97_io_configuration),
    .io_inputs_5(Multiplexer_97_io_inputs_5),
    .io_inputs_4(Multiplexer_97_io_inputs_4),
    .io_inputs_3(Multiplexer_97_io_inputs_3),
    .io_inputs_2(Multiplexer_97_io_inputs_2),
    .io_inputs_1(Multiplexer_97_io_inputs_1),
    .io_inputs_0(Multiplexer_97_io_inputs_0),
    .io_outs_0(Multiplexer_97_io_outs_0)
  );
  Multiplexer_8 Multiplexer_98 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_98_io_configuration),
    .io_inputs_5(Multiplexer_98_io_inputs_5),
    .io_inputs_4(Multiplexer_98_io_inputs_4),
    .io_inputs_3(Multiplexer_98_io_inputs_3),
    .io_inputs_2(Multiplexer_98_io_inputs_2),
    .io_inputs_1(Multiplexer_98_io_inputs_1),
    .io_inputs_0(Multiplexer_98_io_inputs_0),
    .io_outs_0(Multiplexer_98_io_outs_0)
  );
  Multiplexer_8 Multiplexer_99 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_99_io_configuration),
    .io_inputs_5(Multiplexer_99_io_inputs_5),
    .io_inputs_4(Multiplexer_99_io_inputs_4),
    .io_inputs_3(Multiplexer_99_io_inputs_3),
    .io_inputs_2(Multiplexer_99_io_inputs_2),
    .io_inputs_1(Multiplexer_99_io_inputs_1),
    .io_inputs_0(Multiplexer_99_io_inputs_0),
    .io_outs_0(Multiplexer_99_io_outs_0)
  );
  Multiplexer_5 Multiplexer_100 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_100_io_configuration),
    .io_inputs_1(Multiplexer_100_io_inputs_1),
    .io_inputs_0(Multiplexer_100_io_inputs_0),
    .io_outs_0(Multiplexer_100_io_outs_0)
  );
  Multiplexer_5 Multiplexer_101 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_101_io_configuration),
    .io_inputs_1(Multiplexer_101_io_inputs_1),
    .io_inputs_0(Multiplexer_101_io_inputs_0),
    .io_outs_0(Multiplexer_101_io_outs_0)
  );
  Multiplexer_5 Multiplexer_102 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_102_io_configuration),
    .io_inputs_1(Multiplexer_102_io_inputs_1),
    .io_inputs_0(Multiplexer_102_io_inputs_0),
    .io_outs_0(Multiplexer_102_io_outs_0)
  );
  Multiplexer_5 Multiplexer_103 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_103_io_configuration),
    .io_inputs_1(Multiplexer_103_io_inputs_1),
    .io_inputs_0(Multiplexer_103_io_inputs_0),
    .io_outs_0(Multiplexer_103_io_outs_0)
  );
  Multiplexer Multiplexer_104 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_104_io_configuration),
    .io_inputs_4(Multiplexer_104_io_inputs_4),
    .io_inputs_3(Multiplexer_104_io_inputs_3),
    .io_inputs_2(Multiplexer_104_io_inputs_2),
    .io_inputs_1(Multiplexer_104_io_inputs_1),
    .io_inputs_0(Multiplexer_104_io_inputs_0),
    .io_outs_0(Multiplexer_104_io_outs_0)
  );
  Multiplexer Multiplexer_105 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_105_io_configuration),
    .io_inputs_4(Multiplexer_105_io_inputs_4),
    .io_inputs_3(Multiplexer_105_io_inputs_3),
    .io_inputs_2(Multiplexer_105_io_inputs_2),
    .io_inputs_1(Multiplexer_105_io_inputs_1),
    .io_inputs_0(Multiplexer_105_io_inputs_0),
    .io_outs_0(Multiplexer_105_io_outs_0)
  );
  Multiplexer Multiplexer_106 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_106_io_configuration),
    .io_inputs_4(Multiplexer_106_io_inputs_4),
    .io_inputs_3(Multiplexer_106_io_inputs_3),
    .io_inputs_2(Multiplexer_106_io_inputs_2),
    .io_inputs_1(Multiplexer_106_io_inputs_1),
    .io_inputs_0(Multiplexer_106_io_inputs_0),
    .io_outs_0(Multiplexer_106_io_outs_0)
  );
  Multiplexer Multiplexer_107 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_107_io_configuration),
    .io_inputs_4(Multiplexer_107_io_inputs_4),
    .io_inputs_3(Multiplexer_107_io_inputs_3),
    .io_inputs_2(Multiplexer_107_io_inputs_2),
    .io_inputs_1(Multiplexer_107_io_inputs_1),
    .io_inputs_0(Multiplexer_107_io_inputs_0),
    .io_outs_0(Multiplexer_107_io_outs_0)
  );
  Multiplexer Multiplexer_108 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_108_io_configuration),
    .io_inputs_4(Multiplexer_108_io_inputs_4),
    .io_inputs_3(Multiplexer_108_io_inputs_3),
    .io_inputs_2(Multiplexer_108_io_inputs_2),
    .io_inputs_1(Multiplexer_108_io_inputs_1),
    .io_inputs_0(Multiplexer_108_io_inputs_0),
    .io_outs_0(Multiplexer_108_io_outs_0)
  );
  Multiplexer_5 Multiplexer_109 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_109_io_configuration),
    .io_inputs_1(Multiplexer_109_io_inputs_1),
    .io_inputs_0(Multiplexer_109_io_inputs_0),
    .io_outs_0(Multiplexer_109_io_outs_0)
  );
  Multiplexer_5 Multiplexer_110 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_110_io_configuration),
    .io_inputs_1(Multiplexer_110_io_inputs_1),
    .io_inputs_0(Multiplexer_110_io_inputs_0),
    .io_outs_0(Multiplexer_110_io_outs_0)
  );
  Multiplexer_5 Multiplexer_111 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_111_io_configuration),
    .io_inputs_1(Multiplexer_111_io_inputs_1),
    .io_inputs_0(Multiplexer_111_io_inputs_0),
    .io_outs_0(Multiplexer_111_io_outs_0)
  );
  Multiplexer Multiplexer_112 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_112_io_configuration),
    .io_inputs_4(Multiplexer_112_io_inputs_4),
    .io_inputs_3(Multiplexer_112_io_inputs_3),
    .io_inputs_2(Multiplexer_112_io_inputs_2),
    .io_inputs_1(Multiplexer_112_io_inputs_1),
    .io_inputs_0(Multiplexer_112_io_inputs_0),
    .io_outs_0(Multiplexer_112_io_outs_0)
  );
  Multiplexer Multiplexer_113 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_113_io_configuration),
    .io_inputs_4(Multiplexer_113_io_inputs_4),
    .io_inputs_3(Multiplexer_113_io_inputs_3),
    .io_inputs_2(Multiplexer_113_io_inputs_2),
    .io_inputs_1(Multiplexer_113_io_inputs_1),
    .io_inputs_0(Multiplexer_113_io_inputs_0),
    .io_outs_0(Multiplexer_113_io_outs_0)
  );
  Multiplexer Multiplexer_114 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_114_io_configuration),
    .io_inputs_4(Multiplexer_114_io_inputs_4),
    .io_inputs_3(Multiplexer_114_io_inputs_3),
    .io_inputs_2(Multiplexer_114_io_inputs_2),
    .io_inputs_1(Multiplexer_114_io_inputs_1),
    .io_inputs_0(Multiplexer_114_io_inputs_0),
    .io_outs_0(Multiplexer_114_io_outs_0)
  );
  Multiplexer Multiplexer_115 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_115_io_configuration),
    .io_inputs_4(Multiplexer_115_io_inputs_4),
    .io_inputs_3(Multiplexer_115_io_inputs_3),
    .io_inputs_2(Multiplexer_115_io_inputs_2),
    .io_inputs_1(Multiplexer_115_io_inputs_1),
    .io_inputs_0(Multiplexer_115_io_inputs_0),
    .io_outs_0(Multiplexer_115_io_outs_0)
  );
  Multiplexer Multiplexer_116 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_116_io_configuration),
    .io_inputs_4(Multiplexer_116_io_inputs_4),
    .io_inputs_3(Multiplexer_116_io_inputs_3),
    .io_inputs_2(Multiplexer_116_io_inputs_2),
    .io_inputs_1(Multiplexer_116_io_inputs_1),
    .io_inputs_0(Multiplexer_116_io_inputs_0),
    .io_outs_0(Multiplexer_116_io_outs_0)
  );
  Multiplexer_5 Multiplexer_117 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_117_io_configuration),
    .io_inputs_1(Multiplexer_117_io_inputs_1),
    .io_inputs_0(Multiplexer_117_io_inputs_0),
    .io_outs_0(Multiplexer_117_io_outs_0)
  );
  Multiplexer_5 Multiplexer_118 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_118_io_configuration),
    .io_inputs_1(Multiplexer_118_io_inputs_1),
    .io_inputs_0(Multiplexer_118_io_inputs_0),
    .io_outs_0(Multiplexer_118_io_outs_0)
  );
  Multiplexer_5 Multiplexer_119 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_119_io_configuration),
    .io_inputs_1(Multiplexer_119_io_inputs_1),
    .io_inputs_0(Multiplexer_119_io_inputs_0),
    .io_outs_0(Multiplexer_119_io_outs_0)
  );
  Multiplexer_8 Multiplexer_120 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_120_io_configuration),
    .io_inputs_5(Multiplexer_120_io_inputs_5),
    .io_inputs_4(Multiplexer_120_io_inputs_4),
    .io_inputs_3(Multiplexer_120_io_inputs_3),
    .io_inputs_2(Multiplexer_120_io_inputs_2),
    .io_inputs_1(Multiplexer_120_io_inputs_1),
    .io_inputs_0(Multiplexer_120_io_inputs_0),
    .io_outs_0(Multiplexer_120_io_outs_0)
  );
  Multiplexer_8 Multiplexer_121 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_121_io_configuration),
    .io_inputs_5(Multiplexer_121_io_inputs_5),
    .io_inputs_4(Multiplexer_121_io_inputs_4),
    .io_inputs_3(Multiplexer_121_io_inputs_3),
    .io_inputs_2(Multiplexer_121_io_inputs_2),
    .io_inputs_1(Multiplexer_121_io_inputs_1),
    .io_inputs_0(Multiplexer_121_io_inputs_0),
    .io_outs_0(Multiplexer_121_io_outs_0)
  );
  Multiplexer_8 Multiplexer_122 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_122_io_configuration),
    .io_inputs_5(Multiplexer_122_io_inputs_5),
    .io_inputs_4(Multiplexer_122_io_inputs_4),
    .io_inputs_3(Multiplexer_122_io_inputs_3),
    .io_inputs_2(Multiplexer_122_io_inputs_2),
    .io_inputs_1(Multiplexer_122_io_inputs_1),
    .io_inputs_0(Multiplexer_122_io_inputs_0),
    .io_outs_0(Multiplexer_122_io_outs_0)
  );
  Multiplexer_8 Multiplexer_123 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_123_io_configuration),
    .io_inputs_5(Multiplexer_123_io_inputs_5),
    .io_inputs_4(Multiplexer_123_io_inputs_4),
    .io_inputs_3(Multiplexer_123_io_inputs_3),
    .io_inputs_2(Multiplexer_123_io_inputs_2),
    .io_inputs_1(Multiplexer_123_io_inputs_1),
    .io_inputs_0(Multiplexer_123_io_inputs_0),
    .io_outs_0(Multiplexer_123_io_outs_0)
  );
  Multiplexer_8 Multiplexer_124 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_124_io_configuration),
    .io_inputs_5(Multiplexer_124_io_inputs_5),
    .io_inputs_4(Multiplexer_124_io_inputs_4),
    .io_inputs_3(Multiplexer_124_io_inputs_3),
    .io_inputs_2(Multiplexer_124_io_inputs_2),
    .io_inputs_1(Multiplexer_124_io_inputs_1),
    .io_inputs_0(Multiplexer_124_io_inputs_0),
    .io_outs_0(Multiplexer_124_io_outs_0)
  );
  Multiplexer_8 Multiplexer_125 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_125_io_configuration),
    .io_inputs_5(Multiplexer_125_io_inputs_5),
    .io_inputs_4(Multiplexer_125_io_inputs_4),
    .io_inputs_3(Multiplexer_125_io_inputs_3),
    .io_inputs_2(Multiplexer_125_io_inputs_2),
    .io_inputs_1(Multiplexer_125_io_inputs_1),
    .io_inputs_0(Multiplexer_125_io_inputs_0),
    .io_outs_0(Multiplexer_125_io_outs_0)
  );
  Multiplexer_5 Multiplexer_126 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_126_io_configuration),
    .io_inputs_1(Multiplexer_126_io_inputs_1),
    .io_inputs_0(Multiplexer_126_io_inputs_0),
    .io_outs_0(Multiplexer_126_io_outs_0)
  );
  Multiplexer_5 Multiplexer_127 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_127_io_configuration),
    .io_inputs_1(Multiplexer_127_io_inputs_1),
    .io_inputs_0(Multiplexer_127_io_inputs_0),
    .io_outs_0(Multiplexer_127_io_outs_0)
  );
  Multiplexer_5 Multiplexer_128 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_128_io_configuration),
    .io_inputs_1(Multiplexer_128_io_inputs_1),
    .io_inputs_0(Multiplexer_128_io_inputs_0),
    .io_outs_0(Multiplexer_128_io_outs_0)
  );
  Multiplexer_5 Multiplexer_129 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_129_io_configuration),
    .io_inputs_1(Multiplexer_129_io_inputs_1),
    .io_inputs_0(Multiplexer_129_io_inputs_0),
    .io_outs_0(Multiplexer_129_io_outs_0)
  );
  Multiplexer_8 Multiplexer_130 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_130_io_configuration),
    .io_inputs_5(Multiplexer_130_io_inputs_5),
    .io_inputs_4(Multiplexer_130_io_inputs_4),
    .io_inputs_3(Multiplexer_130_io_inputs_3),
    .io_inputs_2(Multiplexer_130_io_inputs_2),
    .io_inputs_1(Multiplexer_130_io_inputs_1),
    .io_inputs_0(Multiplexer_130_io_inputs_0),
    .io_outs_0(Multiplexer_130_io_outs_0)
  );
  Multiplexer_8 Multiplexer_131 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_131_io_configuration),
    .io_inputs_5(Multiplexer_131_io_inputs_5),
    .io_inputs_4(Multiplexer_131_io_inputs_4),
    .io_inputs_3(Multiplexer_131_io_inputs_3),
    .io_inputs_2(Multiplexer_131_io_inputs_2),
    .io_inputs_1(Multiplexer_131_io_inputs_1),
    .io_inputs_0(Multiplexer_131_io_inputs_0),
    .io_outs_0(Multiplexer_131_io_outs_0)
  );
  Multiplexer_8 Multiplexer_132 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_132_io_configuration),
    .io_inputs_5(Multiplexer_132_io_inputs_5),
    .io_inputs_4(Multiplexer_132_io_inputs_4),
    .io_inputs_3(Multiplexer_132_io_inputs_3),
    .io_inputs_2(Multiplexer_132_io_inputs_2),
    .io_inputs_1(Multiplexer_132_io_inputs_1),
    .io_inputs_0(Multiplexer_132_io_inputs_0),
    .io_outs_0(Multiplexer_132_io_outs_0)
  );
  Multiplexer_8 Multiplexer_133 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_133_io_configuration),
    .io_inputs_5(Multiplexer_133_io_inputs_5),
    .io_inputs_4(Multiplexer_133_io_inputs_4),
    .io_inputs_3(Multiplexer_133_io_inputs_3),
    .io_inputs_2(Multiplexer_133_io_inputs_2),
    .io_inputs_1(Multiplexer_133_io_inputs_1),
    .io_inputs_0(Multiplexer_133_io_inputs_0),
    .io_outs_0(Multiplexer_133_io_outs_0)
  );
  Multiplexer_8 Multiplexer_134 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_134_io_configuration),
    .io_inputs_5(Multiplexer_134_io_inputs_5),
    .io_inputs_4(Multiplexer_134_io_inputs_4),
    .io_inputs_3(Multiplexer_134_io_inputs_3),
    .io_inputs_2(Multiplexer_134_io_inputs_2),
    .io_inputs_1(Multiplexer_134_io_inputs_1),
    .io_inputs_0(Multiplexer_134_io_inputs_0),
    .io_outs_0(Multiplexer_134_io_outs_0)
  );
  Multiplexer_8 Multiplexer_135 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_135_io_configuration),
    .io_inputs_5(Multiplexer_135_io_inputs_5),
    .io_inputs_4(Multiplexer_135_io_inputs_4),
    .io_inputs_3(Multiplexer_135_io_inputs_3),
    .io_inputs_2(Multiplexer_135_io_inputs_2),
    .io_inputs_1(Multiplexer_135_io_inputs_1),
    .io_inputs_0(Multiplexer_135_io_inputs_0),
    .io_outs_0(Multiplexer_135_io_outs_0)
  );
  Multiplexer_5 Multiplexer_136 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_136_io_configuration),
    .io_inputs_1(Multiplexer_136_io_inputs_1),
    .io_inputs_0(Multiplexer_136_io_inputs_0),
    .io_outs_0(Multiplexer_136_io_outs_0)
  );
  Multiplexer_5 Multiplexer_137 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_137_io_configuration),
    .io_inputs_1(Multiplexer_137_io_inputs_1),
    .io_inputs_0(Multiplexer_137_io_inputs_0),
    .io_outs_0(Multiplexer_137_io_outs_0)
  );
  Multiplexer_5 Multiplexer_138 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_138_io_configuration),
    .io_inputs_1(Multiplexer_138_io_inputs_1),
    .io_inputs_0(Multiplexer_138_io_inputs_0),
    .io_outs_0(Multiplexer_138_io_outs_0)
  );
  Multiplexer_5 Multiplexer_139 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_139_io_configuration),
    .io_inputs_1(Multiplexer_139_io_inputs_1),
    .io_inputs_0(Multiplexer_139_io_inputs_0),
    .io_outs_0(Multiplexer_139_io_outs_0)
  );
  Multiplexer_8 Multiplexer_140 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_140_io_configuration),
    .io_inputs_5(Multiplexer_140_io_inputs_5),
    .io_inputs_4(Multiplexer_140_io_inputs_4),
    .io_inputs_3(Multiplexer_140_io_inputs_3),
    .io_inputs_2(Multiplexer_140_io_inputs_2),
    .io_inputs_1(Multiplexer_140_io_inputs_1),
    .io_inputs_0(Multiplexer_140_io_inputs_0),
    .io_outs_0(Multiplexer_140_io_outs_0)
  );
  Multiplexer_8 Multiplexer_141 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_141_io_configuration),
    .io_inputs_5(Multiplexer_141_io_inputs_5),
    .io_inputs_4(Multiplexer_141_io_inputs_4),
    .io_inputs_3(Multiplexer_141_io_inputs_3),
    .io_inputs_2(Multiplexer_141_io_inputs_2),
    .io_inputs_1(Multiplexer_141_io_inputs_1),
    .io_inputs_0(Multiplexer_141_io_inputs_0),
    .io_outs_0(Multiplexer_141_io_outs_0)
  );
  Multiplexer_8 Multiplexer_142 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_142_io_configuration),
    .io_inputs_5(Multiplexer_142_io_inputs_5),
    .io_inputs_4(Multiplexer_142_io_inputs_4),
    .io_inputs_3(Multiplexer_142_io_inputs_3),
    .io_inputs_2(Multiplexer_142_io_inputs_2),
    .io_inputs_1(Multiplexer_142_io_inputs_1),
    .io_inputs_0(Multiplexer_142_io_inputs_0),
    .io_outs_0(Multiplexer_142_io_outs_0)
  );
  Multiplexer_8 Multiplexer_143 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_143_io_configuration),
    .io_inputs_5(Multiplexer_143_io_inputs_5),
    .io_inputs_4(Multiplexer_143_io_inputs_4),
    .io_inputs_3(Multiplexer_143_io_inputs_3),
    .io_inputs_2(Multiplexer_143_io_inputs_2),
    .io_inputs_1(Multiplexer_143_io_inputs_1),
    .io_inputs_0(Multiplexer_143_io_inputs_0),
    .io_outs_0(Multiplexer_143_io_outs_0)
  );
  Multiplexer_8 Multiplexer_144 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_144_io_configuration),
    .io_inputs_5(Multiplexer_144_io_inputs_5),
    .io_inputs_4(Multiplexer_144_io_inputs_4),
    .io_inputs_3(Multiplexer_144_io_inputs_3),
    .io_inputs_2(Multiplexer_144_io_inputs_2),
    .io_inputs_1(Multiplexer_144_io_inputs_1),
    .io_inputs_0(Multiplexer_144_io_inputs_0),
    .io_outs_0(Multiplexer_144_io_outs_0)
  );
  Multiplexer_8 Multiplexer_145 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_145_io_configuration),
    .io_inputs_5(Multiplexer_145_io_inputs_5),
    .io_inputs_4(Multiplexer_145_io_inputs_4),
    .io_inputs_3(Multiplexer_145_io_inputs_3),
    .io_inputs_2(Multiplexer_145_io_inputs_2),
    .io_inputs_1(Multiplexer_145_io_inputs_1),
    .io_inputs_0(Multiplexer_145_io_inputs_0),
    .io_outs_0(Multiplexer_145_io_outs_0)
  );
  Multiplexer_5 Multiplexer_146 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_146_io_configuration),
    .io_inputs_1(Multiplexer_146_io_inputs_1),
    .io_inputs_0(Multiplexer_146_io_inputs_0),
    .io_outs_0(Multiplexer_146_io_outs_0)
  );
  Multiplexer_5 Multiplexer_147 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_147_io_configuration),
    .io_inputs_1(Multiplexer_147_io_inputs_1),
    .io_inputs_0(Multiplexer_147_io_inputs_0),
    .io_outs_0(Multiplexer_147_io_outs_0)
  );
  Multiplexer_5 Multiplexer_148 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_148_io_configuration),
    .io_inputs_1(Multiplexer_148_io_inputs_1),
    .io_inputs_0(Multiplexer_148_io_inputs_0),
    .io_outs_0(Multiplexer_148_io_outs_0)
  );
  Multiplexer_5 Multiplexer_149 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_149_io_configuration),
    .io_inputs_1(Multiplexer_149_io_inputs_1),
    .io_inputs_0(Multiplexer_149_io_inputs_0),
    .io_outs_0(Multiplexer_149_io_outs_0)
  );
  Multiplexer_8 Multiplexer_150 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_150_io_configuration),
    .io_inputs_5(Multiplexer_150_io_inputs_5),
    .io_inputs_4(Multiplexer_150_io_inputs_4),
    .io_inputs_3(Multiplexer_150_io_inputs_3),
    .io_inputs_2(Multiplexer_150_io_inputs_2),
    .io_inputs_1(Multiplexer_150_io_inputs_1),
    .io_inputs_0(Multiplexer_150_io_inputs_0),
    .io_outs_0(Multiplexer_150_io_outs_0)
  );
  Multiplexer_8 Multiplexer_151 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_151_io_configuration),
    .io_inputs_5(Multiplexer_151_io_inputs_5),
    .io_inputs_4(Multiplexer_151_io_inputs_4),
    .io_inputs_3(Multiplexer_151_io_inputs_3),
    .io_inputs_2(Multiplexer_151_io_inputs_2),
    .io_inputs_1(Multiplexer_151_io_inputs_1),
    .io_inputs_0(Multiplexer_151_io_inputs_0),
    .io_outs_0(Multiplexer_151_io_outs_0)
  );
  Multiplexer_8 Multiplexer_152 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_152_io_configuration),
    .io_inputs_5(Multiplexer_152_io_inputs_5),
    .io_inputs_4(Multiplexer_152_io_inputs_4),
    .io_inputs_3(Multiplexer_152_io_inputs_3),
    .io_inputs_2(Multiplexer_152_io_inputs_2),
    .io_inputs_1(Multiplexer_152_io_inputs_1),
    .io_inputs_0(Multiplexer_152_io_inputs_0),
    .io_outs_0(Multiplexer_152_io_outs_0)
  );
  Multiplexer_8 Multiplexer_153 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_153_io_configuration),
    .io_inputs_5(Multiplexer_153_io_inputs_5),
    .io_inputs_4(Multiplexer_153_io_inputs_4),
    .io_inputs_3(Multiplexer_153_io_inputs_3),
    .io_inputs_2(Multiplexer_153_io_inputs_2),
    .io_inputs_1(Multiplexer_153_io_inputs_1),
    .io_inputs_0(Multiplexer_153_io_inputs_0),
    .io_outs_0(Multiplexer_153_io_outs_0)
  );
  Multiplexer_8 Multiplexer_154 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_154_io_configuration),
    .io_inputs_5(Multiplexer_154_io_inputs_5),
    .io_inputs_4(Multiplexer_154_io_inputs_4),
    .io_inputs_3(Multiplexer_154_io_inputs_3),
    .io_inputs_2(Multiplexer_154_io_inputs_2),
    .io_inputs_1(Multiplexer_154_io_inputs_1),
    .io_inputs_0(Multiplexer_154_io_inputs_0),
    .io_outs_0(Multiplexer_154_io_outs_0)
  );
  Multiplexer_8 Multiplexer_155 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_155_io_configuration),
    .io_inputs_5(Multiplexer_155_io_inputs_5),
    .io_inputs_4(Multiplexer_155_io_inputs_4),
    .io_inputs_3(Multiplexer_155_io_inputs_3),
    .io_inputs_2(Multiplexer_155_io_inputs_2),
    .io_inputs_1(Multiplexer_155_io_inputs_1),
    .io_inputs_0(Multiplexer_155_io_inputs_0),
    .io_outs_0(Multiplexer_155_io_outs_0)
  );
  Multiplexer_5 Multiplexer_156 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_156_io_configuration),
    .io_inputs_1(Multiplexer_156_io_inputs_1),
    .io_inputs_0(Multiplexer_156_io_inputs_0),
    .io_outs_0(Multiplexer_156_io_outs_0)
  );
  Multiplexer_5 Multiplexer_157 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_157_io_configuration),
    .io_inputs_1(Multiplexer_157_io_inputs_1),
    .io_inputs_0(Multiplexer_157_io_inputs_0),
    .io_outs_0(Multiplexer_157_io_outs_0)
  );
  Multiplexer_5 Multiplexer_158 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_158_io_configuration),
    .io_inputs_1(Multiplexer_158_io_inputs_1),
    .io_inputs_0(Multiplexer_158_io_inputs_0),
    .io_outs_0(Multiplexer_158_io_outs_0)
  );
  Multiplexer_5 Multiplexer_159 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_159_io_configuration),
    .io_inputs_1(Multiplexer_159_io_inputs_1),
    .io_inputs_0(Multiplexer_159_io_inputs_0),
    .io_outs_0(Multiplexer_159_io_outs_0)
  );
  Multiplexer Multiplexer_160 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_160_io_configuration),
    .io_inputs_4(Multiplexer_160_io_inputs_4),
    .io_inputs_3(Multiplexer_160_io_inputs_3),
    .io_inputs_2(Multiplexer_160_io_inputs_2),
    .io_inputs_1(Multiplexer_160_io_inputs_1),
    .io_inputs_0(Multiplexer_160_io_inputs_0),
    .io_outs_0(Multiplexer_160_io_outs_0)
  );
  Multiplexer Multiplexer_161 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_161_io_configuration),
    .io_inputs_4(Multiplexer_161_io_inputs_4),
    .io_inputs_3(Multiplexer_161_io_inputs_3),
    .io_inputs_2(Multiplexer_161_io_inputs_2),
    .io_inputs_1(Multiplexer_161_io_inputs_1),
    .io_inputs_0(Multiplexer_161_io_inputs_0),
    .io_outs_0(Multiplexer_161_io_outs_0)
  );
  Multiplexer Multiplexer_162 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_162_io_configuration),
    .io_inputs_4(Multiplexer_162_io_inputs_4),
    .io_inputs_3(Multiplexer_162_io_inputs_3),
    .io_inputs_2(Multiplexer_162_io_inputs_2),
    .io_inputs_1(Multiplexer_162_io_inputs_1),
    .io_inputs_0(Multiplexer_162_io_inputs_0),
    .io_outs_0(Multiplexer_162_io_outs_0)
  );
  Multiplexer Multiplexer_163 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_163_io_configuration),
    .io_inputs_4(Multiplexer_163_io_inputs_4),
    .io_inputs_3(Multiplexer_163_io_inputs_3),
    .io_inputs_2(Multiplexer_163_io_inputs_2),
    .io_inputs_1(Multiplexer_163_io_inputs_1),
    .io_inputs_0(Multiplexer_163_io_inputs_0),
    .io_outs_0(Multiplexer_163_io_outs_0)
  );
  Multiplexer Multiplexer_164 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_164_io_configuration),
    .io_inputs_4(Multiplexer_164_io_inputs_4),
    .io_inputs_3(Multiplexer_164_io_inputs_3),
    .io_inputs_2(Multiplexer_164_io_inputs_2),
    .io_inputs_1(Multiplexer_164_io_inputs_1),
    .io_inputs_0(Multiplexer_164_io_inputs_0),
    .io_outs_0(Multiplexer_164_io_outs_0)
  );
  Multiplexer_5 Multiplexer_165 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_165_io_configuration),
    .io_inputs_1(Multiplexer_165_io_inputs_1),
    .io_inputs_0(Multiplexer_165_io_inputs_0),
    .io_outs_0(Multiplexer_165_io_outs_0)
  );
  Multiplexer_5 Multiplexer_166 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_166_io_configuration),
    .io_inputs_1(Multiplexer_166_io_inputs_1),
    .io_inputs_0(Multiplexer_166_io_inputs_0),
    .io_outs_0(Multiplexer_166_io_outs_0)
  );
  Multiplexer_5 Multiplexer_167 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_167_io_configuration),
    .io_inputs_1(Multiplexer_167_io_inputs_1),
    .io_inputs_0(Multiplexer_167_io_inputs_0),
    .io_outs_0(Multiplexer_167_io_outs_0)
  );
  Multiplexer Multiplexer_168 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_168_io_configuration),
    .io_inputs_4(Multiplexer_168_io_inputs_4),
    .io_inputs_3(Multiplexer_168_io_inputs_3),
    .io_inputs_2(Multiplexer_168_io_inputs_2),
    .io_inputs_1(Multiplexer_168_io_inputs_1),
    .io_inputs_0(Multiplexer_168_io_inputs_0),
    .io_outs_0(Multiplexer_168_io_outs_0)
  );
  Multiplexer Multiplexer_169 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_169_io_configuration),
    .io_inputs_4(Multiplexer_169_io_inputs_4),
    .io_inputs_3(Multiplexer_169_io_inputs_3),
    .io_inputs_2(Multiplexer_169_io_inputs_2),
    .io_inputs_1(Multiplexer_169_io_inputs_1),
    .io_inputs_0(Multiplexer_169_io_inputs_0),
    .io_outs_0(Multiplexer_169_io_outs_0)
  );
  Multiplexer Multiplexer_170 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_170_io_configuration),
    .io_inputs_4(Multiplexer_170_io_inputs_4),
    .io_inputs_3(Multiplexer_170_io_inputs_3),
    .io_inputs_2(Multiplexer_170_io_inputs_2),
    .io_inputs_1(Multiplexer_170_io_inputs_1),
    .io_inputs_0(Multiplexer_170_io_inputs_0),
    .io_outs_0(Multiplexer_170_io_outs_0)
  );
  Multiplexer Multiplexer_171 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_171_io_configuration),
    .io_inputs_4(Multiplexer_171_io_inputs_4),
    .io_inputs_3(Multiplexer_171_io_inputs_3),
    .io_inputs_2(Multiplexer_171_io_inputs_2),
    .io_inputs_1(Multiplexer_171_io_inputs_1),
    .io_inputs_0(Multiplexer_171_io_inputs_0),
    .io_outs_0(Multiplexer_171_io_outs_0)
  );
  Multiplexer Multiplexer_172 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_172_io_configuration),
    .io_inputs_4(Multiplexer_172_io_inputs_4),
    .io_inputs_3(Multiplexer_172_io_inputs_3),
    .io_inputs_2(Multiplexer_172_io_inputs_2),
    .io_inputs_1(Multiplexer_172_io_inputs_1),
    .io_inputs_0(Multiplexer_172_io_inputs_0),
    .io_outs_0(Multiplexer_172_io_outs_0)
  );
  Multiplexer_5 Multiplexer_173 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_173_io_configuration),
    .io_inputs_1(Multiplexer_173_io_inputs_1),
    .io_inputs_0(Multiplexer_173_io_inputs_0),
    .io_outs_0(Multiplexer_173_io_outs_0)
  );
  Multiplexer_5 Multiplexer_174 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_174_io_configuration),
    .io_inputs_1(Multiplexer_174_io_inputs_1),
    .io_inputs_0(Multiplexer_174_io_inputs_0),
    .io_outs_0(Multiplexer_174_io_outs_0)
  );
  Multiplexer_5 Multiplexer_175 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_175_io_configuration),
    .io_inputs_1(Multiplexer_175_io_inputs_1),
    .io_inputs_0(Multiplexer_175_io_inputs_0),
    .io_outs_0(Multiplexer_175_io_outs_0)
  );
  Multiplexer_8 Multiplexer_176 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_176_io_configuration),
    .io_inputs_5(Multiplexer_176_io_inputs_5),
    .io_inputs_4(Multiplexer_176_io_inputs_4),
    .io_inputs_3(Multiplexer_176_io_inputs_3),
    .io_inputs_2(Multiplexer_176_io_inputs_2),
    .io_inputs_1(Multiplexer_176_io_inputs_1),
    .io_inputs_0(Multiplexer_176_io_inputs_0),
    .io_outs_0(Multiplexer_176_io_outs_0)
  );
  Multiplexer_8 Multiplexer_177 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_177_io_configuration),
    .io_inputs_5(Multiplexer_177_io_inputs_5),
    .io_inputs_4(Multiplexer_177_io_inputs_4),
    .io_inputs_3(Multiplexer_177_io_inputs_3),
    .io_inputs_2(Multiplexer_177_io_inputs_2),
    .io_inputs_1(Multiplexer_177_io_inputs_1),
    .io_inputs_0(Multiplexer_177_io_inputs_0),
    .io_outs_0(Multiplexer_177_io_outs_0)
  );
  Multiplexer_8 Multiplexer_178 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_178_io_configuration),
    .io_inputs_5(Multiplexer_178_io_inputs_5),
    .io_inputs_4(Multiplexer_178_io_inputs_4),
    .io_inputs_3(Multiplexer_178_io_inputs_3),
    .io_inputs_2(Multiplexer_178_io_inputs_2),
    .io_inputs_1(Multiplexer_178_io_inputs_1),
    .io_inputs_0(Multiplexer_178_io_inputs_0),
    .io_outs_0(Multiplexer_178_io_outs_0)
  );
  Multiplexer_8 Multiplexer_179 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_179_io_configuration),
    .io_inputs_5(Multiplexer_179_io_inputs_5),
    .io_inputs_4(Multiplexer_179_io_inputs_4),
    .io_inputs_3(Multiplexer_179_io_inputs_3),
    .io_inputs_2(Multiplexer_179_io_inputs_2),
    .io_inputs_1(Multiplexer_179_io_inputs_1),
    .io_inputs_0(Multiplexer_179_io_inputs_0),
    .io_outs_0(Multiplexer_179_io_outs_0)
  );
  Multiplexer_8 Multiplexer_180 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_180_io_configuration),
    .io_inputs_5(Multiplexer_180_io_inputs_5),
    .io_inputs_4(Multiplexer_180_io_inputs_4),
    .io_inputs_3(Multiplexer_180_io_inputs_3),
    .io_inputs_2(Multiplexer_180_io_inputs_2),
    .io_inputs_1(Multiplexer_180_io_inputs_1),
    .io_inputs_0(Multiplexer_180_io_inputs_0),
    .io_outs_0(Multiplexer_180_io_outs_0)
  );
  Multiplexer_8 Multiplexer_181 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_181_io_configuration),
    .io_inputs_5(Multiplexer_181_io_inputs_5),
    .io_inputs_4(Multiplexer_181_io_inputs_4),
    .io_inputs_3(Multiplexer_181_io_inputs_3),
    .io_inputs_2(Multiplexer_181_io_inputs_2),
    .io_inputs_1(Multiplexer_181_io_inputs_1),
    .io_inputs_0(Multiplexer_181_io_inputs_0),
    .io_outs_0(Multiplexer_181_io_outs_0)
  );
  Multiplexer_5 Multiplexer_182 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_182_io_configuration),
    .io_inputs_1(Multiplexer_182_io_inputs_1),
    .io_inputs_0(Multiplexer_182_io_inputs_0),
    .io_outs_0(Multiplexer_182_io_outs_0)
  );
  Multiplexer_5 Multiplexer_183 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_183_io_configuration),
    .io_inputs_1(Multiplexer_183_io_inputs_1),
    .io_inputs_0(Multiplexer_183_io_inputs_0),
    .io_outs_0(Multiplexer_183_io_outs_0)
  );
  Multiplexer_5 Multiplexer_184 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_184_io_configuration),
    .io_inputs_1(Multiplexer_184_io_inputs_1),
    .io_inputs_0(Multiplexer_184_io_inputs_0),
    .io_outs_0(Multiplexer_184_io_outs_0)
  );
  Multiplexer_5 Multiplexer_185 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_185_io_configuration),
    .io_inputs_1(Multiplexer_185_io_inputs_1),
    .io_inputs_0(Multiplexer_185_io_inputs_0),
    .io_outs_0(Multiplexer_185_io_outs_0)
  );
  Multiplexer_8 Multiplexer_186 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_186_io_configuration),
    .io_inputs_5(Multiplexer_186_io_inputs_5),
    .io_inputs_4(Multiplexer_186_io_inputs_4),
    .io_inputs_3(Multiplexer_186_io_inputs_3),
    .io_inputs_2(Multiplexer_186_io_inputs_2),
    .io_inputs_1(Multiplexer_186_io_inputs_1),
    .io_inputs_0(Multiplexer_186_io_inputs_0),
    .io_outs_0(Multiplexer_186_io_outs_0)
  );
  Multiplexer_8 Multiplexer_187 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_187_io_configuration),
    .io_inputs_5(Multiplexer_187_io_inputs_5),
    .io_inputs_4(Multiplexer_187_io_inputs_4),
    .io_inputs_3(Multiplexer_187_io_inputs_3),
    .io_inputs_2(Multiplexer_187_io_inputs_2),
    .io_inputs_1(Multiplexer_187_io_inputs_1),
    .io_inputs_0(Multiplexer_187_io_inputs_0),
    .io_outs_0(Multiplexer_187_io_outs_0)
  );
  Multiplexer_8 Multiplexer_188 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_188_io_configuration),
    .io_inputs_5(Multiplexer_188_io_inputs_5),
    .io_inputs_4(Multiplexer_188_io_inputs_4),
    .io_inputs_3(Multiplexer_188_io_inputs_3),
    .io_inputs_2(Multiplexer_188_io_inputs_2),
    .io_inputs_1(Multiplexer_188_io_inputs_1),
    .io_inputs_0(Multiplexer_188_io_inputs_0),
    .io_outs_0(Multiplexer_188_io_outs_0)
  );
  Multiplexer_8 Multiplexer_189 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_189_io_configuration),
    .io_inputs_5(Multiplexer_189_io_inputs_5),
    .io_inputs_4(Multiplexer_189_io_inputs_4),
    .io_inputs_3(Multiplexer_189_io_inputs_3),
    .io_inputs_2(Multiplexer_189_io_inputs_2),
    .io_inputs_1(Multiplexer_189_io_inputs_1),
    .io_inputs_0(Multiplexer_189_io_inputs_0),
    .io_outs_0(Multiplexer_189_io_outs_0)
  );
  Multiplexer_8 Multiplexer_190 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_190_io_configuration),
    .io_inputs_5(Multiplexer_190_io_inputs_5),
    .io_inputs_4(Multiplexer_190_io_inputs_4),
    .io_inputs_3(Multiplexer_190_io_inputs_3),
    .io_inputs_2(Multiplexer_190_io_inputs_2),
    .io_inputs_1(Multiplexer_190_io_inputs_1),
    .io_inputs_0(Multiplexer_190_io_inputs_0),
    .io_outs_0(Multiplexer_190_io_outs_0)
  );
  Multiplexer_8 Multiplexer_191 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_191_io_configuration),
    .io_inputs_5(Multiplexer_191_io_inputs_5),
    .io_inputs_4(Multiplexer_191_io_inputs_4),
    .io_inputs_3(Multiplexer_191_io_inputs_3),
    .io_inputs_2(Multiplexer_191_io_inputs_2),
    .io_inputs_1(Multiplexer_191_io_inputs_1),
    .io_inputs_0(Multiplexer_191_io_inputs_0),
    .io_outs_0(Multiplexer_191_io_outs_0)
  );
  Multiplexer_5 Multiplexer_192 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_192_io_configuration),
    .io_inputs_1(Multiplexer_192_io_inputs_1),
    .io_inputs_0(Multiplexer_192_io_inputs_0),
    .io_outs_0(Multiplexer_192_io_outs_0)
  );
  Multiplexer_5 Multiplexer_193 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_193_io_configuration),
    .io_inputs_1(Multiplexer_193_io_inputs_1),
    .io_inputs_0(Multiplexer_193_io_inputs_0),
    .io_outs_0(Multiplexer_193_io_outs_0)
  );
  Multiplexer_5 Multiplexer_194 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_194_io_configuration),
    .io_inputs_1(Multiplexer_194_io_inputs_1),
    .io_inputs_0(Multiplexer_194_io_inputs_0),
    .io_outs_0(Multiplexer_194_io_outs_0)
  );
  Multiplexer_5 Multiplexer_195 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_195_io_configuration),
    .io_inputs_1(Multiplexer_195_io_inputs_1),
    .io_inputs_0(Multiplexer_195_io_inputs_0),
    .io_outs_0(Multiplexer_195_io_outs_0)
  );
  Multiplexer_8 Multiplexer_196 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_196_io_configuration),
    .io_inputs_5(Multiplexer_196_io_inputs_5),
    .io_inputs_4(Multiplexer_196_io_inputs_4),
    .io_inputs_3(Multiplexer_196_io_inputs_3),
    .io_inputs_2(Multiplexer_196_io_inputs_2),
    .io_inputs_1(Multiplexer_196_io_inputs_1),
    .io_inputs_0(Multiplexer_196_io_inputs_0),
    .io_outs_0(Multiplexer_196_io_outs_0)
  );
  Multiplexer_8 Multiplexer_197 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_197_io_configuration),
    .io_inputs_5(Multiplexer_197_io_inputs_5),
    .io_inputs_4(Multiplexer_197_io_inputs_4),
    .io_inputs_3(Multiplexer_197_io_inputs_3),
    .io_inputs_2(Multiplexer_197_io_inputs_2),
    .io_inputs_1(Multiplexer_197_io_inputs_1),
    .io_inputs_0(Multiplexer_197_io_inputs_0),
    .io_outs_0(Multiplexer_197_io_outs_0)
  );
  Multiplexer_8 Multiplexer_198 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_198_io_configuration),
    .io_inputs_5(Multiplexer_198_io_inputs_5),
    .io_inputs_4(Multiplexer_198_io_inputs_4),
    .io_inputs_3(Multiplexer_198_io_inputs_3),
    .io_inputs_2(Multiplexer_198_io_inputs_2),
    .io_inputs_1(Multiplexer_198_io_inputs_1),
    .io_inputs_0(Multiplexer_198_io_inputs_0),
    .io_outs_0(Multiplexer_198_io_outs_0)
  );
  Multiplexer_8 Multiplexer_199 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_199_io_configuration),
    .io_inputs_5(Multiplexer_199_io_inputs_5),
    .io_inputs_4(Multiplexer_199_io_inputs_4),
    .io_inputs_3(Multiplexer_199_io_inputs_3),
    .io_inputs_2(Multiplexer_199_io_inputs_2),
    .io_inputs_1(Multiplexer_199_io_inputs_1),
    .io_inputs_0(Multiplexer_199_io_inputs_0),
    .io_outs_0(Multiplexer_199_io_outs_0)
  );
  Multiplexer_8 Multiplexer_200 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_200_io_configuration),
    .io_inputs_5(Multiplexer_200_io_inputs_5),
    .io_inputs_4(Multiplexer_200_io_inputs_4),
    .io_inputs_3(Multiplexer_200_io_inputs_3),
    .io_inputs_2(Multiplexer_200_io_inputs_2),
    .io_inputs_1(Multiplexer_200_io_inputs_1),
    .io_inputs_0(Multiplexer_200_io_inputs_0),
    .io_outs_0(Multiplexer_200_io_outs_0)
  );
  Multiplexer_8 Multiplexer_201 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_201_io_configuration),
    .io_inputs_5(Multiplexer_201_io_inputs_5),
    .io_inputs_4(Multiplexer_201_io_inputs_4),
    .io_inputs_3(Multiplexer_201_io_inputs_3),
    .io_inputs_2(Multiplexer_201_io_inputs_2),
    .io_inputs_1(Multiplexer_201_io_inputs_1),
    .io_inputs_0(Multiplexer_201_io_inputs_0),
    .io_outs_0(Multiplexer_201_io_outs_0)
  );
  Multiplexer_5 Multiplexer_202 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_202_io_configuration),
    .io_inputs_1(Multiplexer_202_io_inputs_1),
    .io_inputs_0(Multiplexer_202_io_inputs_0),
    .io_outs_0(Multiplexer_202_io_outs_0)
  );
  Multiplexer_5 Multiplexer_203 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_203_io_configuration),
    .io_inputs_1(Multiplexer_203_io_inputs_1),
    .io_inputs_0(Multiplexer_203_io_inputs_0),
    .io_outs_0(Multiplexer_203_io_outs_0)
  );
  Multiplexer_5 Multiplexer_204 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_204_io_configuration),
    .io_inputs_1(Multiplexer_204_io_inputs_1),
    .io_inputs_0(Multiplexer_204_io_inputs_0),
    .io_outs_0(Multiplexer_204_io_outs_0)
  );
  Multiplexer_5 Multiplexer_205 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_205_io_configuration),
    .io_inputs_1(Multiplexer_205_io_inputs_1),
    .io_inputs_0(Multiplexer_205_io_inputs_0),
    .io_outs_0(Multiplexer_205_io_outs_0)
  );
  Multiplexer_8 Multiplexer_206 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_206_io_configuration),
    .io_inputs_5(Multiplexer_206_io_inputs_5),
    .io_inputs_4(Multiplexer_206_io_inputs_4),
    .io_inputs_3(Multiplexer_206_io_inputs_3),
    .io_inputs_2(Multiplexer_206_io_inputs_2),
    .io_inputs_1(Multiplexer_206_io_inputs_1),
    .io_inputs_0(Multiplexer_206_io_inputs_0),
    .io_outs_0(Multiplexer_206_io_outs_0)
  );
  Multiplexer_8 Multiplexer_207 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_207_io_configuration),
    .io_inputs_5(Multiplexer_207_io_inputs_5),
    .io_inputs_4(Multiplexer_207_io_inputs_4),
    .io_inputs_3(Multiplexer_207_io_inputs_3),
    .io_inputs_2(Multiplexer_207_io_inputs_2),
    .io_inputs_1(Multiplexer_207_io_inputs_1),
    .io_inputs_0(Multiplexer_207_io_inputs_0),
    .io_outs_0(Multiplexer_207_io_outs_0)
  );
  Multiplexer_8 Multiplexer_208 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_208_io_configuration),
    .io_inputs_5(Multiplexer_208_io_inputs_5),
    .io_inputs_4(Multiplexer_208_io_inputs_4),
    .io_inputs_3(Multiplexer_208_io_inputs_3),
    .io_inputs_2(Multiplexer_208_io_inputs_2),
    .io_inputs_1(Multiplexer_208_io_inputs_1),
    .io_inputs_0(Multiplexer_208_io_inputs_0),
    .io_outs_0(Multiplexer_208_io_outs_0)
  );
  Multiplexer_8 Multiplexer_209 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_209_io_configuration),
    .io_inputs_5(Multiplexer_209_io_inputs_5),
    .io_inputs_4(Multiplexer_209_io_inputs_4),
    .io_inputs_3(Multiplexer_209_io_inputs_3),
    .io_inputs_2(Multiplexer_209_io_inputs_2),
    .io_inputs_1(Multiplexer_209_io_inputs_1),
    .io_inputs_0(Multiplexer_209_io_inputs_0),
    .io_outs_0(Multiplexer_209_io_outs_0)
  );
  Multiplexer_8 Multiplexer_210 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_210_io_configuration),
    .io_inputs_5(Multiplexer_210_io_inputs_5),
    .io_inputs_4(Multiplexer_210_io_inputs_4),
    .io_inputs_3(Multiplexer_210_io_inputs_3),
    .io_inputs_2(Multiplexer_210_io_inputs_2),
    .io_inputs_1(Multiplexer_210_io_inputs_1),
    .io_inputs_0(Multiplexer_210_io_inputs_0),
    .io_outs_0(Multiplexer_210_io_outs_0)
  );
  Multiplexer_8 Multiplexer_211 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_211_io_configuration),
    .io_inputs_5(Multiplexer_211_io_inputs_5),
    .io_inputs_4(Multiplexer_211_io_inputs_4),
    .io_inputs_3(Multiplexer_211_io_inputs_3),
    .io_inputs_2(Multiplexer_211_io_inputs_2),
    .io_inputs_1(Multiplexer_211_io_inputs_1),
    .io_inputs_0(Multiplexer_211_io_inputs_0),
    .io_outs_0(Multiplexer_211_io_outs_0)
  );
  Multiplexer_5 Multiplexer_212 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_212_io_configuration),
    .io_inputs_1(Multiplexer_212_io_inputs_1),
    .io_inputs_0(Multiplexer_212_io_inputs_0),
    .io_outs_0(Multiplexer_212_io_outs_0)
  );
  Multiplexer_5 Multiplexer_213 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_213_io_configuration),
    .io_inputs_1(Multiplexer_213_io_inputs_1),
    .io_inputs_0(Multiplexer_213_io_inputs_0),
    .io_outs_0(Multiplexer_213_io_outs_0)
  );
  Multiplexer_5 Multiplexer_214 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_214_io_configuration),
    .io_inputs_1(Multiplexer_214_io_inputs_1),
    .io_inputs_0(Multiplexer_214_io_inputs_0),
    .io_outs_0(Multiplexer_214_io_outs_0)
  );
  Multiplexer_5 Multiplexer_215 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_215_io_configuration),
    .io_inputs_1(Multiplexer_215_io_inputs_1),
    .io_inputs_0(Multiplexer_215_io_inputs_0),
    .io_outs_0(Multiplexer_215_io_outs_0)
  );
  Multiplexer Multiplexer_216 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_216_io_configuration),
    .io_inputs_4(Multiplexer_216_io_inputs_4),
    .io_inputs_3(Multiplexer_216_io_inputs_3),
    .io_inputs_2(Multiplexer_216_io_inputs_2),
    .io_inputs_1(Multiplexer_216_io_inputs_1),
    .io_inputs_0(Multiplexer_216_io_inputs_0),
    .io_outs_0(Multiplexer_216_io_outs_0)
  );
  Multiplexer Multiplexer_217 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_217_io_configuration),
    .io_inputs_4(Multiplexer_217_io_inputs_4),
    .io_inputs_3(Multiplexer_217_io_inputs_3),
    .io_inputs_2(Multiplexer_217_io_inputs_2),
    .io_inputs_1(Multiplexer_217_io_inputs_1),
    .io_inputs_0(Multiplexer_217_io_inputs_0),
    .io_outs_0(Multiplexer_217_io_outs_0)
  );
  Multiplexer Multiplexer_218 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_218_io_configuration),
    .io_inputs_4(Multiplexer_218_io_inputs_4),
    .io_inputs_3(Multiplexer_218_io_inputs_3),
    .io_inputs_2(Multiplexer_218_io_inputs_2),
    .io_inputs_1(Multiplexer_218_io_inputs_1),
    .io_inputs_0(Multiplexer_218_io_inputs_0),
    .io_outs_0(Multiplexer_218_io_outs_0)
  );
  Multiplexer Multiplexer_219 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_219_io_configuration),
    .io_inputs_4(Multiplexer_219_io_inputs_4),
    .io_inputs_3(Multiplexer_219_io_inputs_3),
    .io_inputs_2(Multiplexer_219_io_inputs_2),
    .io_inputs_1(Multiplexer_219_io_inputs_1),
    .io_inputs_0(Multiplexer_219_io_inputs_0),
    .io_outs_0(Multiplexer_219_io_outs_0)
  );
  Multiplexer Multiplexer_220 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_220_io_configuration),
    .io_inputs_4(Multiplexer_220_io_inputs_4),
    .io_inputs_3(Multiplexer_220_io_inputs_3),
    .io_inputs_2(Multiplexer_220_io_inputs_2),
    .io_inputs_1(Multiplexer_220_io_inputs_1),
    .io_inputs_0(Multiplexer_220_io_inputs_0),
    .io_outs_0(Multiplexer_220_io_outs_0)
  );
  Multiplexer_5 Multiplexer_221 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_221_io_configuration),
    .io_inputs_1(Multiplexer_221_io_inputs_1),
    .io_inputs_0(Multiplexer_221_io_inputs_0),
    .io_outs_0(Multiplexer_221_io_outs_0)
  );
  Multiplexer_5 Multiplexer_222 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_222_io_configuration),
    .io_inputs_1(Multiplexer_222_io_inputs_1),
    .io_inputs_0(Multiplexer_222_io_inputs_0),
    .io_outs_0(Multiplexer_222_io_outs_0)
  );
  Multiplexer_5 Multiplexer_223 ( // @[TopModule.scala 169:11]
    .io_configuration(Multiplexer_223_io_configuration),
    .io_inputs_1(Multiplexer_223_io_inputs_1),
    .io_inputs_0(Multiplexer_223_io_inputs_0),
    .io_outs_0(Multiplexer_223_io_outs_0)
  );
  ConstUnit ConstUnit ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_io_configuration),
    .io_outs_0(ConstUnit_io_outs_0)
  );
  ConstUnit ConstUnit_1 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_1_io_configuration),
    .io_outs_0(ConstUnit_1_io_outs_0)
  );
  ConstUnit ConstUnit_2 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_2_io_configuration),
    .io_outs_0(ConstUnit_2_io_outs_0)
  );
  ConstUnit ConstUnit_3 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_3_io_configuration),
    .io_outs_0(ConstUnit_3_io_outs_0)
  );
  ConstUnit ConstUnit_4 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_4_io_configuration),
    .io_outs_0(ConstUnit_4_io_outs_0)
  );
  ConstUnit ConstUnit_5 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_5_io_configuration),
    .io_outs_0(ConstUnit_5_io_outs_0)
  );
  ConstUnit ConstUnit_6 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_6_io_configuration),
    .io_outs_0(ConstUnit_6_io_outs_0)
  );
  ConstUnit ConstUnit_7 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_7_io_configuration),
    .io_outs_0(ConstUnit_7_io_outs_0)
  );
  ConstUnit ConstUnit_8 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_8_io_configuration),
    .io_outs_0(ConstUnit_8_io_outs_0)
  );
  ConstUnit ConstUnit_9 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_9_io_configuration),
    .io_outs_0(ConstUnit_9_io_outs_0)
  );
  ConstUnit ConstUnit_10 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_10_io_configuration),
    .io_outs_0(ConstUnit_10_io_outs_0)
  );
  ConstUnit ConstUnit_11 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_11_io_configuration),
    .io_outs_0(ConstUnit_11_io_outs_0)
  );
  ConstUnit ConstUnit_12 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_12_io_configuration),
    .io_outs_0(ConstUnit_12_io_outs_0)
  );
  ConstUnit ConstUnit_13 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_13_io_configuration),
    .io_outs_0(ConstUnit_13_io_outs_0)
  );
  ConstUnit ConstUnit_14 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_14_io_configuration),
    .io_outs_0(ConstUnit_14_io_outs_0)
  );
  ConstUnit ConstUnit_15 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_15_io_configuration),
    .io_outs_0(ConstUnit_15_io_outs_0)
  );
  ConstUnit ConstUnit_16 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_16_io_configuration),
    .io_outs_0(ConstUnit_16_io_outs_0)
  );
  ConstUnit ConstUnit_17 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_17_io_configuration),
    .io_outs_0(ConstUnit_17_io_outs_0)
  );
  ConstUnit ConstUnit_18 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_18_io_configuration),
    .io_outs_0(ConstUnit_18_io_outs_0)
  );
  ConstUnit ConstUnit_19 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_19_io_configuration),
    .io_outs_0(ConstUnit_19_io_outs_0)
  );
  ConstUnit ConstUnit_20 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_20_io_configuration),
    .io_outs_0(ConstUnit_20_io_outs_0)
  );
  ConstUnit ConstUnit_21 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_21_io_configuration),
    .io_outs_0(ConstUnit_21_io_outs_0)
  );
  ConstUnit ConstUnit_22 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_22_io_configuration),
    .io_outs_0(ConstUnit_22_io_outs_0)
  );
  ConstUnit ConstUnit_23 ( // @[TopModule.scala 177:21]
    .io_configuration(ConstUnit_23_io_configuration),
    .io_outs_0(ConstUnit_23_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_clock),
    .reset(LoadStoreUnit_reset),
    .io_configuration(LoadStoreUnit_io_configuration),
    .io_en(LoadStoreUnit_io_en),
    .io_skewing(LoadStoreUnit_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_io_streamIn_bits),
    .io_len(LoadStoreUnit_io_len),
    .io_streamOut_ready(LoadStoreUnit_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_io_streamOut_bits),
    .io_base(LoadStoreUnit_io_base),
    .io_start(LoadStoreUnit_io_start),
    .io_enqEn(LoadStoreUnit_io_enqEn),
    .io_deqEn(LoadStoreUnit_io_deqEn),
    .io_idle(LoadStoreUnit_io_idle),
    .io_inputs_1(LoadStoreUnit_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_io_inputs_0),
    .io_outs_0(LoadStoreUnit_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_1 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_1_clock),
    .reset(LoadStoreUnit_1_reset),
    .io_configuration(LoadStoreUnit_1_io_configuration),
    .io_en(LoadStoreUnit_1_io_en),
    .io_skewing(LoadStoreUnit_1_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_1_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_1_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_1_io_streamIn_bits),
    .io_len(LoadStoreUnit_1_io_len),
    .io_streamOut_ready(LoadStoreUnit_1_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_1_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_1_io_streamOut_bits),
    .io_base(LoadStoreUnit_1_io_base),
    .io_start(LoadStoreUnit_1_io_start),
    .io_enqEn(LoadStoreUnit_1_io_enqEn),
    .io_deqEn(LoadStoreUnit_1_io_deqEn),
    .io_idle(LoadStoreUnit_1_io_idle),
    .io_inputs_1(LoadStoreUnit_1_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_1_io_inputs_0),
    .io_outs_0(LoadStoreUnit_1_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_2 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_2_clock),
    .reset(LoadStoreUnit_2_reset),
    .io_configuration(LoadStoreUnit_2_io_configuration),
    .io_en(LoadStoreUnit_2_io_en),
    .io_skewing(LoadStoreUnit_2_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_2_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_2_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_2_io_streamIn_bits),
    .io_len(LoadStoreUnit_2_io_len),
    .io_streamOut_ready(LoadStoreUnit_2_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_2_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_2_io_streamOut_bits),
    .io_base(LoadStoreUnit_2_io_base),
    .io_start(LoadStoreUnit_2_io_start),
    .io_enqEn(LoadStoreUnit_2_io_enqEn),
    .io_deqEn(LoadStoreUnit_2_io_deqEn),
    .io_idle(LoadStoreUnit_2_io_idle),
    .io_inputs_1(LoadStoreUnit_2_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_2_io_inputs_0),
    .io_outs_0(LoadStoreUnit_2_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_3 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_3_clock),
    .reset(LoadStoreUnit_3_reset),
    .io_configuration(LoadStoreUnit_3_io_configuration),
    .io_en(LoadStoreUnit_3_io_en),
    .io_skewing(LoadStoreUnit_3_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_3_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_3_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_3_io_streamIn_bits),
    .io_len(LoadStoreUnit_3_io_len),
    .io_streamOut_ready(LoadStoreUnit_3_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_3_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_3_io_streamOut_bits),
    .io_base(LoadStoreUnit_3_io_base),
    .io_start(LoadStoreUnit_3_io_start),
    .io_enqEn(LoadStoreUnit_3_io_enqEn),
    .io_deqEn(LoadStoreUnit_3_io_deqEn),
    .io_idle(LoadStoreUnit_3_io_idle),
    .io_inputs_1(LoadStoreUnit_3_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_3_io_inputs_0),
    .io_outs_0(LoadStoreUnit_3_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_4 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_4_clock),
    .reset(LoadStoreUnit_4_reset),
    .io_configuration(LoadStoreUnit_4_io_configuration),
    .io_en(LoadStoreUnit_4_io_en),
    .io_skewing(LoadStoreUnit_4_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_4_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_4_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_4_io_streamIn_bits),
    .io_len(LoadStoreUnit_4_io_len),
    .io_streamOut_ready(LoadStoreUnit_4_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_4_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_4_io_streamOut_bits),
    .io_base(LoadStoreUnit_4_io_base),
    .io_start(LoadStoreUnit_4_io_start),
    .io_enqEn(LoadStoreUnit_4_io_enqEn),
    .io_deqEn(LoadStoreUnit_4_io_deqEn),
    .io_idle(LoadStoreUnit_4_io_idle),
    .io_inputs_1(LoadStoreUnit_4_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_4_io_inputs_0),
    .io_outs_0(LoadStoreUnit_4_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_5 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_5_clock),
    .reset(LoadStoreUnit_5_reset),
    .io_configuration(LoadStoreUnit_5_io_configuration),
    .io_en(LoadStoreUnit_5_io_en),
    .io_skewing(LoadStoreUnit_5_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_5_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_5_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_5_io_streamIn_bits),
    .io_len(LoadStoreUnit_5_io_len),
    .io_streamOut_ready(LoadStoreUnit_5_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_5_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_5_io_streamOut_bits),
    .io_base(LoadStoreUnit_5_io_base),
    .io_start(LoadStoreUnit_5_io_start),
    .io_enqEn(LoadStoreUnit_5_io_enqEn),
    .io_deqEn(LoadStoreUnit_5_io_deqEn),
    .io_idle(LoadStoreUnit_5_io_idle),
    .io_inputs_1(LoadStoreUnit_5_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_5_io_inputs_0),
    .io_outs_0(LoadStoreUnit_5_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_6 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_6_clock),
    .reset(LoadStoreUnit_6_reset),
    .io_configuration(LoadStoreUnit_6_io_configuration),
    .io_en(LoadStoreUnit_6_io_en),
    .io_skewing(LoadStoreUnit_6_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_6_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_6_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_6_io_streamIn_bits),
    .io_len(LoadStoreUnit_6_io_len),
    .io_streamOut_ready(LoadStoreUnit_6_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_6_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_6_io_streamOut_bits),
    .io_base(LoadStoreUnit_6_io_base),
    .io_start(LoadStoreUnit_6_io_start),
    .io_enqEn(LoadStoreUnit_6_io_enqEn),
    .io_deqEn(LoadStoreUnit_6_io_deqEn),
    .io_idle(LoadStoreUnit_6_io_idle),
    .io_inputs_1(LoadStoreUnit_6_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_6_io_inputs_0),
    .io_outs_0(LoadStoreUnit_6_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_7 ( // @[TopModule.scala 186:21]
    .clock(LoadStoreUnit_7_clock),
    .reset(LoadStoreUnit_7_reset),
    .io_configuration(LoadStoreUnit_7_io_configuration),
    .io_en(LoadStoreUnit_7_io_en),
    .io_skewing(LoadStoreUnit_7_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_7_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_7_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_7_io_streamIn_bits),
    .io_len(LoadStoreUnit_7_io_len),
    .io_streamOut_ready(LoadStoreUnit_7_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_7_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_7_io_streamOut_bits),
    .io_base(LoadStoreUnit_7_io_base),
    .io_start(LoadStoreUnit_7_io_start),
    .io_enqEn(LoadStoreUnit_7_io_enqEn),
    .io_deqEn(LoadStoreUnit_7_io_deqEn),
    .io_idle(LoadStoreUnit_7_io_idle),
    .io_inputs_1(LoadStoreUnit_7_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_7_io_inputs_0),
    .io_outs_0(LoadStoreUnit_7_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController_16 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_16_clock),
    .reset(MultiIIScheduleController_16_reset),
    .io_en(MultiIIScheduleController_16_io_en),
    .io_schedules_0(MultiIIScheduleController_16_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_16_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_16_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_16_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_16_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_16_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_16_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_16_io_schedules_7),
    .io_II(MultiIIScheduleController_16_io_II),
    .io_valid(MultiIIScheduleController_16_io_valid),
    .io_skewing(MultiIIScheduleController_16_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_17 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_17_clock),
    .reset(MultiIIScheduleController_17_reset),
    .io_en(MultiIIScheduleController_17_io_en),
    .io_schedules_0(MultiIIScheduleController_17_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_17_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_17_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_17_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_17_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_17_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_17_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_17_io_schedules_7),
    .io_II(MultiIIScheduleController_17_io_II),
    .io_valid(MultiIIScheduleController_17_io_valid),
    .io_skewing(MultiIIScheduleController_17_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_18 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_18_clock),
    .reset(MultiIIScheduleController_18_reset),
    .io_en(MultiIIScheduleController_18_io_en),
    .io_schedules_0(MultiIIScheduleController_18_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_18_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_18_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_18_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_18_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_18_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_18_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_18_io_schedules_7),
    .io_II(MultiIIScheduleController_18_io_II),
    .io_valid(MultiIIScheduleController_18_io_valid),
    .io_skewing(MultiIIScheduleController_18_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_19 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_19_clock),
    .reset(MultiIIScheduleController_19_reset),
    .io_en(MultiIIScheduleController_19_io_en),
    .io_schedules_0(MultiIIScheduleController_19_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_19_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_19_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_19_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_19_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_19_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_19_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_19_io_schedules_7),
    .io_II(MultiIIScheduleController_19_io_II),
    .io_valid(MultiIIScheduleController_19_io_valid),
    .io_skewing(MultiIIScheduleController_19_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_20 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_20_clock),
    .reset(MultiIIScheduleController_20_reset),
    .io_en(MultiIIScheduleController_20_io_en),
    .io_schedules_0(MultiIIScheduleController_20_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_20_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_20_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_20_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_20_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_20_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_20_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_20_io_schedules_7),
    .io_II(MultiIIScheduleController_20_io_II),
    .io_valid(MultiIIScheduleController_20_io_valid),
    .io_skewing(MultiIIScheduleController_20_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_21 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_21_clock),
    .reset(MultiIIScheduleController_21_reset),
    .io_en(MultiIIScheduleController_21_io_en),
    .io_schedules_0(MultiIIScheduleController_21_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_21_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_21_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_21_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_21_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_21_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_21_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_21_io_schedules_7),
    .io_II(MultiIIScheduleController_21_io_II),
    .io_valid(MultiIIScheduleController_21_io_valid),
    .io_skewing(MultiIIScheduleController_21_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_22 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_22_clock),
    .reset(MultiIIScheduleController_22_reset),
    .io_en(MultiIIScheduleController_22_io_en),
    .io_schedules_0(MultiIIScheduleController_22_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_22_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_22_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_22_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_22_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_22_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_22_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_22_io_schedules_7),
    .io_II(MultiIIScheduleController_22_io_II),
    .io_valid(MultiIIScheduleController_22_io_valid),
    .io_skewing(MultiIIScheduleController_22_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_23 ( // @[TopModule.scala 200:23]
    .clock(MultiIIScheduleController_23_clock),
    .reset(MultiIIScheduleController_23_reset),
    .io_en(MultiIIScheduleController_23_io_en),
    .io_schedules_0(MultiIIScheduleController_23_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_23_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_23_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_23_io_schedules_3),
    .io_schedules_4(MultiIIScheduleController_23_io_schedules_4),
    .io_schedules_5(MultiIIScheduleController_23_io_schedules_5),
    .io_schedules_6(MultiIIScheduleController_23_io_schedules_6),
    .io_schedules_7(MultiIIScheduleController_23_io_schedules_7),
    .io_II(MultiIIScheduleController_23_io_II),
    .io_valid(MultiIIScheduleController_23_io_valid),
    .io_skewing(MultiIIScheduleController_23_io_skewing)
  );
  ConfigController configControllers_0 ( // @[TopModule.scala 262:34]
    .clock(configControllers_0_clock),
    .reset(configControllers_0_reset),
    .io_en(configControllers_0_io_en),
    .io_II(configControllers_0_io_II),
    .io_inConfig(configControllers_0_io_inConfig),
    .io_outConfig(configControllers_0_io_outConfig)
  );
  Dispatch_145 Dispatch_1 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_1_io_configuration),
    .io_outs_11(Dispatch_1_io_outs_11),
    .io_outs_10(Dispatch_1_io_outs_10),
    .io_outs_9(Dispatch_1_io_outs_9),
    .io_outs_8(Dispatch_1_io_outs_8),
    .io_outs_7(Dispatch_1_io_outs_7),
    .io_outs_6(Dispatch_1_io_outs_6),
    .io_outs_5(Dispatch_1_io_outs_5),
    .io_outs_4(Dispatch_1_io_outs_4),
    .io_outs_3(Dispatch_1_io_outs_3),
    .io_outs_2(Dispatch_1_io_outs_2),
    .io_outs_1(Dispatch_1_io_outs_1),
    .io_outs_0(Dispatch_1_io_outs_0)
  );
  ConfigController configControllers_1 ( // @[TopModule.scala 262:34]
    .clock(configControllers_1_clock),
    .reset(configControllers_1_reset),
    .io_en(configControllers_1_io_en),
    .io_II(configControllers_1_io_II),
    .io_inConfig(configControllers_1_io_inConfig),
    .io_outConfig(configControllers_1_io_outConfig)
  );
  Dispatch_145 Dispatch_2 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_2_io_configuration),
    .io_outs_11(Dispatch_2_io_outs_11),
    .io_outs_10(Dispatch_2_io_outs_10),
    .io_outs_9(Dispatch_2_io_outs_9),
    .io_outs_8(Dispatch_2_io_outs_8),
    .io_outs_7(Dispatch_2_io_outs_7),
    .io_outs_6(Dispatch_2_io_outs_6),
    .io_outs_5(Dispatch_2_io_outs_5),
    .io_outs_4(Dispatch_2_io_outs_4),
    .io_outs_3(Dispatch_2_io_outs_3),
    .io_outs_2(Dispatch_2_io_outs_2),
    .io_outs_1(Dispatch_2_io_outs_1),
    .io_outs_0(Dispatch_2_io_outs_0)
  );
  ConfigController_2 configControllers_2 ( // @[TopModule.scala 262:34]
    .clock(configControllers_2_clock),
    .reset(configControllers_2_reset),
    .io_en(configControllers_2_io_en),
    .io_II(configControllers_2_io_II),
    .io_inConfig(configControllers_2_io_inConfig),
    .io_outConfig(configControllers_2_io_outConfig)
  );
  Dispatch_147 Dispatch_3 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_3_io_configuration),
    .io_outs_12(Dispatch_3_io_outs_12),
    .io_outs_11(Dispatch_3_io_outs_11),
    .io_outs_10(Dispatch_3_io_outs_10),
    .io_outs_9(Dispatch_3_io_outs_9),
    .io_outs_8(Dispatch_3_io_outs_8),
    .io_outs_7(Dispatch_3_io_outs_7),
    .io_outs_6(Dispatch_3_io_outs_6),
    .io_outs_5(Dispatch_3_io_outs_5),
    .io_outs_4(Dispatch_3_io_outs_4),
    .io_outs_3(Dispatch_3_io_outs_3),
    .io_outs_2(Dispatch_3_io_outs_2),
    .io_outs_1(Dispatch_3_io_outs_1),
    .io_outs_0(Dispatch_3_io_outs_0)
  );
  ConfigController_3 configControllers_3 ( // @[TopModule.scala 262:34]
    .clock(configControllers_3_clock),
    .reset(configControllers_3_reset),
    .io_en(configControllers_3_io_en),
    .io_II(configControllers_3_io_II),
    .io_inConfig(configControllers_3_io_inConfig),
    .io_outConfig(configControllers_3_io_outConfig)
  );
  Dispatch_148 Dispatch_4 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_4_io_configuration),
    .io_outs_17(Dispatch_4_io_outs_17),
    .io_outs_16(Dispatch_4_io_outs_16),
    .io_outs_15(Dispatch_4_io_outs_15),
    .io_outs_14(Dispatch_4_io_outs_14),
    .io_outs_13(Dispatch_4_io_outs_13),
    .io_outs_12(Dispatch_4_io_outs_12),
    .io_outs_11(Dispatch_4_io_outs_11),
    .io_outs_10(Dispatch_4_io_outs_10),
    .io_outs_9(Dispatch_4_io_outs_9),
    .io_outs_8(Dispatch_4_io_outs_8),
    .io_outs_7(Dispatch_4_io_outs_7),
    .io_outs_6(Dispatch_4_io_outs_6),
    .io_outs_5(Dispatch_4_io_outs_5),
    .io_outs_4(Dispatch_4_io_outs_4),
    .io_outs_3(Dispatch_4_io_outs_3),
    .io_outs_2(Dispatch_4_io_outs_2),
    .io_outs_1(Dispatch_4_io_outs_1),
    .io_outs_0(Dispatch_4_io_outs_0)
  );
  ConfigController_3 configControllers_4 ( // @[TopModule.scala 262:34]
    .clock(configControllers_4_clock),
    .reset(configControllers_4_reset),
    .io_en(configControllers_4_io_en),
    .io_II(configControllers_4_io_II),
    .io_inConfig(configControllers_4_io_inConfig),
    .io_outConfig(configControllers_4_io_outConfig)
  );
  Dispatch_148 Dispatch_5 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_5_io_configuration),
    .io_outs_17(Dispatch_5_io_outs_17),
    .io_outs_16(Dispatch_5_io_outs_16),
    .io_outs_15(Dispatch_5_io_outs_15),
    .io_outs_14(Dispatch_5_io_outs_14),
    .io_outs_13(Dispatch_5_io_outs_13),
    .io_outs_12(Dispatch_5_io_outs_12),
    .io_outs_11(Dispatch_5_io_outs_11),
    .io_outs_10(Dispatch_5_io_outs_10),
    .io_outs_9(Dispatch_5_io_outs_9),
    .io_outs_8(Dispatch_5_io_outs_8),
    .io_outs_7(Dispatch_5_io_outs_7),
    .io_outs_6(Dispatch_5_io_outs_6),
    .io_outs_5(Dispatch_5_io_outs_5),
    .io_outs_4(Dispatch_5_io_outs_4),
    .io_outs_3(Dispatch_5_io_outs_3),
    .io_outs_2(Dispatch_5_io_outs_2),
    .io_outs_1(Dispatch_5_io_outs_1),
    .io_outs_0(Dispatch_5_io_outs_0)
  );
  ConfigController_3 configControllers_5 ( // @[TopModule.scala 262:34]
    .clock(configControllers_5_clock),
    .reset(configControllers_5_reset),
    .io_en(configControllers_5_io_en),
    .io_II(configControllers_5_io_II),
    .io_inConfig(configControllers_5_io_inConfig),
    .io_outConfig(configControllers_5_io_outConfig)
  );
  Dispatch_148 Dispatch_6 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_6_io_configuration),
    .io_outs_17(Dispatch_6_io_outs_17),
    .io_outs_16(Dispatch_6_io_outs_16),
    .io_outs_15(Dispatch_6_io_outs_15),
    .io_outs_14(Dispatch_6_io_outs_14),
    .io_outs_13(Dispatch_6_io_outs_13),
    .io_outs_12(Dispatch_6_io_outs_12),
    .io_outs_11(Dispatch_6_io_outs_11),
    .io_outs_10(Dispatch_6_io_outs_10),
    .io_outs_9(Dispatch_6_io_outs_9),
    .io_outs_8(Dispatch_6_io_outs_8),
    .io_outs_7(Dispatch_6_io_outs_7),
    .io_outs_6(Dispatch_6_io_outs_6),
    .io_outs_5(Dispatch_6_io_outs_5),
    .io_outs_4(Dispatch_6_io_outs_4),
    .io_outs_3(Dispatch_6_io_outs_3),
    .io_outs_2(Dispatch_6_io_outs_2),
    .io_outs_1(Dispatch_6_io_outs_1),
    .io_outs_0(Dispatch_6_io_outs_0)
  );
  ConfigController_3 configControllers_6 ( // @[TopModule.scala 262:34]
    .clock(configControllers_6_clock),
    .reset(configControllers_6_reset),
    .io_en(configControllers_6_io_en),
    .io_II(configControllers_6_io_II),
    .io_inConfig(configControllers_6_io_inConfig),
    .io_outConfig(configControllers_6_io_outConfig)
  );
  Dispatch_148 Dispatch_7 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_7_io_configuration),
    .io_outs_17(Dispatch_7_io_outs_17),
    .io_outs_16(Dispatch_7_io_outs_16),
    .io_outs_15(Dispatch_7_io_outs_15),
    .io_outs_14(Dispatch_7_io_outs_14),
    .io_outs_13(Dispatch_7_io_outs_13),
    .io_outs_12(Dispatch_7_io_outs_12),
    .io_outs_11(Dispatch_7_io_outs_11),
    .io_outs_10(Dispatch_7_io_outs_10),
    .io_outs_9(Dispatch_7_io_outs_9),
    .io_outs_8(Dispatch_7_io_outs_8),
    .io_outs_7(Dispatch_7_io_outs_7),
    .io_outs_6(Dispatch_7_io_outs_6),
    .io_outs_5(Dispatch_7_io_outs_5),
    .io_outs_4(Dispatch_7_io_outs_4),
    .io_outs_3(Dispatch_7_io_outs_3),
    .io_outs_2(Dispatch_7_io_outs_2),
    .io_outs_1(Dispatch_7_io_outs_1),
    .io_outs_0(Dispatch_7_io_outs_0)
  );
  ConfigController_2 configControllers_7 ( // @[TopModule.scala 262:34]
    .clock(configControllers_7_clock),
    .reset(configControllers_7_reset),
    .io_en(configControllers_7_io_en),
    .io_II(configControllers_7_io_II),
    .io_inConfig(configControllers_7_io_inConfig),
    .io_outConfig(configControllers_7_io_outConfig)
  );
  Dispatch_147 Dispatch_8 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_8_io_configuration),
    .io_outs_12(Dispatch_8_io_outs_12),
    .io_outs_11(Dispatch_8_io_outs_11),
    .io_outs_10(Dispatch_8_io_outs_10),
    .io_outs_9(Dispatch_8_io_outs_9),
    .io_outs_8(Dispatch_8_io_outs_8),
    .io_outs_7(Dispatch_8_io_outs_7),
    .io_outs_6(Dispatch_8_io_outs_6),
    .io_outs_5(Dispatch_8_io_outs_5),
    .io_outs_4(Dispatch_8_io_outs_4),
    .io_outs_3(Dispatch_8_io_outs_3),
    .io_outs_2(Dispatch_8_io_outs_2),
    .io_outs_1(Dispatch_8_io_outs_1),
    .io_outs_0(Dispatch_8_io_outs_0)
  );
  ConfigController_2 configControllers_8 ( // @[TopModule.scala 262:34]
    .clock(configControllers_8_clock),
    .reset(configControllers_8_reset),
    .io_en(configControllers_8_io_en),
    .io_II(configControllers_8_io_II),
    .io_inConfig(configControllers_8_io_inConfig),
    .io_outConfig(configControllers_8_io_outConfig)
  );
  Dispatch_147 Dispatch_9 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_9_io_configuration),
    .io_outs_12(Dispatch_9_io_outs_12),
    .io_outs_11(Dispatch_9_io_outs_11),
    .io_outs_10(Dispatch_9_io_outs_10),
    .io_outs_9(Dispatch_9_io_outs_9),
    .io_outs_8(Dispatch_9_io_outs_8),
    .io_outs_7(Dispatch_9_io_outs_7),
    .io_outs_6(Dispatch_9_io_outs_6),
    .io_outs_5(Dispatch_9_io_outs_5),
    .io_outs_4(Dispatch_9_io_outs_4),
    .io_outs_3(Dispatch_9_io_outs_3),
    .io_outs_2(Dispatch_9_io_outs_2),
    .io_outs_1(Dispatch_9_io_outs_1),
    .io_outs_0(Dispatch_9_io_outs_0)
  );
  ConfigController_3 configControllers_9 ( // @[TopModule.scala 262:34]
    .clock(configControllers_9_clock),
    .reset(configControllers_9_reset),
    .io_en(configControllers_9_io_en),
    .io_II(configControllers_9_io_II),
    .io_inConfig(configControllers_9_io_inConfig),
    .io_outConfig(configControllers_9_io_outConfig)
  );
  Dispatch_148 Dispatch_10 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_10_io_configuration),
    .io_outs_17(Dispatch_10_io_outs_17),
    .io_outs_16(Dispatch_10_io_outs_16),
    .io_outs_15(Dispatch_10_io_outs_15),
    .io_outs_14(Dispatch_10_io_outs_14),
    .io_outs_13(Dispatch_10_io_outs_13),
    .io_outs_12(Dispatch_10_io_outs_12),
    .io_outs_11(Dispatch_10_io_outs_11),
    .io_outs_10(Dispatch_10_io_outs_10),
    .io_outs_9(Dispatch_10_io_outs_9),
    .io_outs_8(Dispatch_10_io_outs_8),
    .io_outs_7(Dispatch_10_io_outs_7),
    .io_outs_6(Dispatch_10_io_outs_6),
    .io_outs_5(Dispatch_10_io_outs_5),
    .io_outs_4(Dispatch_10_io_outs_4),
    .io_outs_3(Dispatch_10_io_outs_3),
    .io_outs_2(Dispatch_10_io_outs_2),
    .io_outs_1(Dispatch_10_io_outs_1),
    .io_outs_0(Dispatch_10_io_outs_0)
  );
  ConfigController_3 configControllers_10 ( // @[TopModule.scala 262:34]
    .clock(configControllers_10_clock),
    .reset(configControllers_10_reset),
    .io_en(configControllers_10_io_en),
    .io_II(configControllers_10_io_II),
    .io_inConfig(configControllers_10_io_inConfig),
    .io_outConfig(configControllers_10_io_outConfig)
  );
  Dispatch_148 Dispatch_11 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_11_io_configuration),
    .io_outs_17(Dispatch_11_io_outs_17),
    .io_outs_16(Dispatch_11_io_outs_16),
    .io_outs_15(Dispatch_11_io_outs_15),
    .io_outs_14(Dispatch_11_io_outs_14),
    .io_outs_13(Dispatch_11_io_outs_13),
    .io_outs_12(Dispatch_11_io_outs_12),
    .io_outs_11(Dispatch_11_io_outs_11),
    .io_outs_10(Dispatch_11_io_outs_10),
    .io_outs_9(Dispatch_11_io_outs_9),
    .io_outs_8(Dispatch_11_io_outs_8),
    .io_outs_7(Dispatch_11_io_outs_7),
    .io_outs_6(Dispatch_11_io_outs_6),
    .io_outs_5(Dispatch_11_io_outs_5),
    .io_outs_4(Dispatch_11_io_outs_4),
    .io_outs_3(Dispatch_11_io_outs_3),
    .io_outs_2(Dispatch_11_io_outs_2),
    .io_outs_1(Dispatch_11_io_outs_1),
    .io_outs_0(Dispatch_11_io_outs_0)
  );
  ConfigController_3 configControllers_11 ( // @[TopModule.scala 262:34]
    .clock(configControllers_11_clock),
    .reset(configControllers_11_reset),
    .io_en(configControllers_11_io_en),
    .io_II(configControllers_11_io_II),
    .io_inConfig(configControllers_11_io_inConfig),
    .io_outConfig(configControllers_11_io_outConfig)
  );
  Dispatch_148 Dispatch_12 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_12_io_configuration),
    .io_outs_17(Dispatch_12_io_outs_17),
    .io_outs_16(Dispatch_12_io_outs_16),
    .io_outs_15(Dispatch_12_io_outs_15),
    .io_outs_14(Dispatch_12_io_outs_14),
    .io_outs_13(Dispatch_12_io_outs_13),
    .io_outs_12(Dispatch_12_io_outs_12),
    .io_outs_11(Dispatch_12_io_outs_11),
    .io_outs_10(Dispatch_12_io_outs_10),
    .io_outs_9(Dispatch_12_io_outs_9),
    .io_outs_8(Dispatch_12_io_outs_8),
    .io_outs_7(Dispatch_12_io_outs_7),
    .io_outs_6(Dispatch_12_io_outs_6),
    .io_outs_5(Dispatch_12_io_outs_5),
    .io_outs_4(Dispatch_12_io_outs_4),
    .io_outs_3(Dispatch_12_io_outs_3),
    .io_outs_2(Dispatch_12_io_outs_2),
    .io_outs_1(Dispatch_12_io_outs_1),
    .io_outs_0(Dispatch_12_io_outs_0)
  );
  ConfigController_3 configControllers_12 ( // @[TopModule.scala 262:34]
    .clock(configControllers_12_clock),
    .reset(configControllers_12_reset),
    .io_en(configControllers_12_io_en),
    .io_II(configControllers_12_io_II),
    .io_inConfig(configControllers_12_io_inConfig),
    .io_outConfig(configControllers_12_io_outConfig)
  );
  Dispatch_148 Dispatch_13 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_13_io_configuration),
    .io_outs_17(Dispatch_13_io_outs_17),
    .io_outs_16(Dispatch_13_io_outs_16),
    .io_outs_15(Dispatch_13_io_outs_15),
    .io_outs_14(Dispatch_13_io_outs_14),
    .io_outs_13(Dispatch_13_io_outs_13),
    .io_outs_12(Dispatch_13_io_outs_12),
    .io_outs_11(Dispatch_13_io_outs_11),
    .io_outs_10(Dispatch_13_io_outs_10),
    .io_outs_9(Dispatch_13_io_outs_9),
    .io_outs_8(Dispatch_13_io_outs_8),
    .io_outs_7(Dispatch_13_io_outs_7),
    .io_outs_6(Dispatch_13_io_outs_6),
    .io_outs_5(Dispatch_13_io_outs_5),
    .io_outs_4(Dispatch_13_io_outs_4),
    .io_outs_3(Dispatch_13_io_outs_3),
    .io_outs_2(Dispatch_13_io_outs_2),
    .io_outs_1(Dispatch_13_io_outs_1),
    .io_outs_0(Dispatch_13_io_outs_0)
  );
  ConfigController_2 configControllers_13 ( // @[TopModule.scala 262:34]
    .clock(configControllers_13_clock),
    .reset(configControllers_13_reset),
    .io_en(configControllers_13_io_en),
    .io_II(configControllers_13_io_II),
    .io_inConfig(configControllers_13_io_inConfig),
    .io_outConfig(configControllers_13_io_outConfig)
  );
  Dispatch_147 Dispatch_14 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_14_io_configuration),
    .io_outs_12(Dispatch_14_io_outs_12),
    .io_outs_11(Dispatch_14_io_outs_11),
    .io_outs_10(Dispatch_14_io_outs_10),
    .io_outs_9(Dispatch_14_io_outs_9),
    .io_outs_8(Dispatch_14_io_outs_8),
    .io_outs_7(Dispatch_14_io_outs_7),
    .io_outs_6(Dispatch_14_io_outs_6),
    .io_outs_5(Dispatch_14_io_outs_5),
    .io_outs_4(Dispatch_14_io_outs_4),
    .io_outs_3(Dispatch_14_io_outs_3),
    .io_outs_2(Dispatch_14_io_outs_2),
    .io_outs_1(Dispatch_14_io_outs_1),
    .io_outs_0(Dispatch_14_io_outs_0)
  );
  ConfigController_2 configControllers_14 ( // @[TopModule.scala 262:34]
    .clock(configControllers_14_clock),
    .reset(configControllers_14_reset),
    .io_en(configControllers_14_io_en),
    .io_II(configControllers_14_io_II),
    .io_inConfig(configControllers_14_io_inConfig),
    .io_outConfig(configControllers_14_io_outConfig)
  );
  Dispatch_147 Dispatch_15 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_15_io_configuration),
    .io_outs_12(Dispatch_15_io_outs_12),
    .io_outs_11(Dispatch_15_io_outs_11),
    .io_outs_10(Dispatch_15_io_outs_10),
    .io_outs_9(Dispatch_15_io_outs_9),
    .io_outs_8(Dispatch_15_io_outs_8),
    .io_outs_7(Dispatch_15_io_outs_7),
    .io_outs_6(Dispatch_15_io_outs_6),
    .io_outs_5(Dispatch_15_io_outs_5),
    .io_outs_4(Dispatch_15_io_outs_4),
    .io_outs_3(Dispatch_15_io_outs_3),
    .io_outs_2(Dispatch_15_io_outs_2),
    .io_outs_1(Dispatch_15_io_outs_1),
    .io_outs_0(Dispatch_15_io_outs_0)
  );
  ConfigController_3 configControllers_15 ( // @[TopModule.scala 262:34]
    .clock(configControllers_15_clock),
    .reset(configControllers_15_reset),
    .io_en(configControllers_15_io_en),
    .io_II(configControllers_15_io_II),
    .io_inConfig(configControllers_15_io_inConfig),
    .io_outConfig(configControllers_15_io_outConfig)
  );
  Dispatch_148 Dispatch_16 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_16_io_configuration),
    .io_outs_17(Dispatch_16_io_outs_17),
    .io_outs_16(Dispatch_16_io_outs_16),
    .io_outs_15(Dispatch_16_io_outs_15),
    .io_outs_14(Dispatch_16_io_outs_14),
    .io_outs_13(Dispatch_16_io_outs_13),
    .io_outs_12(Dispatch_16_io_outs_12),
    .io_outs_11(Dispatch_16_io_outs_11),
    .io_outs_10(Dispatch_16_io_outs_10),
    .io_outs_9(Dispatch_16_io_outs_9),
    .io_outs_8(Dispatch_16_io_outs_8),
    .io_outs_7(Dispatch_16_io_outs_7),
    .io_outs_6(Dispatch_16_io_outs_6),
    .io_outs_5(Dispatch_16_io_outs_5),
    .io_outs_4(Dispatch_16_io_outs_4),
    .io_outs_3(Dispatch_16_io_outs_3),
    .io_outs_2(Dispatch_16_io_outs_2),
    .io_outs_1(Dispatch_16_io_outs_1),
    .io_outs_0(Dispatch_16_io_outs_0)
  );
  ConfigController_3 configControllers_16 ( // @[TopModule.scala 262:34]
    .clock(configControllers_16_clock),
    .reset(configControllers_16_reset),
    .io_en(configControllers_16_io_en),
    .io_II(configControllers_16_io_II),
    .io_inConfig(configControllers_16_io_inConfig),
    .io_outConfig(configControllers_16_io_outConfig)
  );
  Dispatch_148 Dispatch_17 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_17_io_configuration),
    .io_outs_17(Dispatch_17_io_outs_17),
    .io_outs_16(Dispatch_17_io_outs_16),
    .io_outs_15(Dispatch_17_io_outs_15),
    .io_outs_14(Dispatch_17_io_outs_14),
    .io_outs_13(Dispatch_17_io_outs_13),
    .io_outs_12(Dispatch_17_io_outs_12),
    .io_outs_11(Dispatch_17_io_outs_11),
    .io_outs_10(Dispatch_17_io_outs_10),
    .io_outs_9(Dispatch_17_io_outs_9),
    .io_outs_8(Dispatch_17_io_outs_8),
    .io_outs_7(Dispatch_17_io_outs_7),
    .io_outs_6(Dispatch_17_io_outs_6),
    .io_outs_5(Dispatch_17_io_outs_5),
    .io_outs_4(Dispatch_17_io_outs_4),
    .io_outs_3(Dispatch_17_io_outs_3),
    .io_outs_2(Dispatch_17_io_outs_2),
    .io_outs_1(Dispatch_17_io_outs_1),
    .io_outs_0(Dispatch_17_io_outs_0)
  );
  ConfigController_3 configControllers_17 ( // @[TopModule.scala 262:34]
    .clock(configControllers_17_clock),
    .reset(configControllers_17_reset),
    .io_en(configControllers_17_io_en),
    .io_II(configControllers_17_io_II),
    .io_inConfig(configControllers_17_io_inConfig),
    .io_outConfig(configControllers_17_io_outConfig)
  );
  Dispatch_148 Dispatch_18 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_18_io_configuration),
    .io_outs_17(Dispatch_18_io_outs_17),
    .io_outs_16(Dispatch_18_io_outs_16),
    .io_outs_15(Dispatch_18_io_outs_15),
    .io_outs_14(Dispatch_18_io_outs_14),
    .io_outs_13(Dispatch_18_io_outs_13),
    .io_outs_12(Dispatch_18_io_outs_12),
    .io_outs_11(Dispatch_18_io_outs_11),
    .io_outs_10(Dispatch_18_io_outs_10),
    .io_outs_9(Dispatch_18_io_outs_9),
    .io_outs_8(Dispatch_18_io_outs_8),
    .io_outs_7(Dispatch_18_io_outs_7),
    .io_outs_6(Dispatch_18_io_outs_6),
    .io_outs_5(Dispatch_18_io_outs_5),
    .io_outs_4(Dispatch_18_io_outs_4),
    .io_outs_3(Dispatch_18_io_outs_3),
    .io_outs_2(Dispatch_18_io_outs_2),
    .io_outs_1(Dispatch_18_io_outs_1),
    .io_outs_0(Dispatch_18_io_outs_0)
  );
  ConfigController_3 configControllers_18 ( // @[TopModule.scala 262:34]
    .clock(configControllers_18_clock),
    .reset(configControllers_18_reset),
    .io_en(configControllers_18_io_en),
    .io_II(configControllers_18_io_II),
    .io_inConfig(configControllers_18_io_inConfig),
    .io_outConfig(configControllers_18_io_outConfig)
  );
  Dispatch_148 Dispatch_19 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_19_io_configuration),
    .io_outs_17(Dispatch_19_io_outs_17),
    .io_outs_16(Dispatch_19_io_outs_16),
    .io_outs_15(Dispatch_19_io_outs_15),
    .io_outs_14(Dispatch_19_io_outs_14),
    .io_outs_13(Dispatch_19_io_outs_13),
    .io_outs_12(Dispatch_19_io_outs_12),
    .io_outs_11(Dispatch_19_io_outs_11),
    .io_outs_10(Dispatch_19_io_outs_10),
    .io_outs_9(Dispatch_19_io_outs_9),
    .io_outs_8(Dispatch_19_io_outs_8),
    .io_outs_7(Dispatch_19_io_outs_7),
    .io_outs_6(Dispatch_19_io_outs_6),
    .io_outs_5(Dispatch_19_io_outs_5),
    .io_outs_4(Dispatch_19_io_outs_4),
    .io_outs_3(Dispatch_19_io_outs_3),
    .io_outs_2(Dispatch_19_io_outs_2),
    .io_outs_1(Dispatch_19_io_outs_1),
    .io_outs_0(Dispatch_19_io_outs_0)
  );
  ConfigController_2 configControllers_19 ( // @[TopModule.scala 262:34]
    .clock(configControllers_19_clock),
    .reset(configControllers_19_reset),
    .io_en(configControllers_19_io_en),
    .io_II(configControllers_19_io_II),
    .io_inConfig(configControllers_19_io_inConfig),
    .io_outConfig(configControllers_19_io_outConfig)
  );
  Dispatch_147 Dispatch_20 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_20_io_configuration),
    .io_outs_12(Dispatch_20_io_outs_12),
    .io_outs_11(Dispatch_20_io_outs_11),
    .io_outs_10(Dispatch_20_io_outs_10),
    .io_outs_9(Dispatch_20_io_outs_9),
    .io_outs_8(Dispatch_20_io_outs_8),
    .io_outs_7(Dispatch_20_io_outs_7),
    .io_outs_6(Dispatch_20_io_outs_6),
    .io_outs_5(Dispatch_20_io_outs_5),
    .io_outs_4(Dispatch_20_io_outs_4),
    .io_outs_3(Dispatch_20_io_outs_3),
    .io_outs_2(Dispatch_20_io_outs_2),
    .io_outs_1(Dispatch_20_io_outs_1),
    .io_outs_0(Dispatch_20_io_outs_0)
  );
  ConfigController_2 configControllers_20 ( // @[TopModule.scala 262:34]
    .clock(configControllers_20_clock),
    .reset(configControllers_20_reset),
    .io_en(configControllers_20_io_en),
    .io_II(configControllers_20_io_II),
    .io_inConfig(configControllers_20_io_inConfig),
    .io_outConfig(configControllers_20_io_outConfig)
  );
  Dispatch_147 Dispatch_21 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_21_io_configuration),
    .io_outs_12(Dispatch_21_io_outs_12),
    .io_outs_11(Dispatch_21_io_outs_11),
    .io_outs_10(Dispatch_21_io_outs_10),
    .io_outs_9(Dispatch_21_io_outs_9),
    .io_outs_8(Dispatch_21_io_outs_8),
    .io_outs_7(Dispatch_21_io_outs_7),
    .io_outs_6(Dispatch_21_io_outs_6),
    .io_outs_5(Dispatch_21_io_outs_5),
    .io_outs_4(Dispatch_21_io_outs_4),
    .io_outs_3(Dispatch_21_io_outs_3),
    .io_outs_2(Dispatch_21_io_outs_2),
    .io_outs_1(Dispatch_21_io_outs_1),
    .io_outs_0(Dispatch_21_io_outs_0)
  );
  ConfigController_3 configControllers_21 ( // @[TopModule.scala 262:34]
    .clock(configControllers_21_clock),
    .reset(configControllers_21_reset),
    .io_en(configControllers_21_io_en),
    .io_II(configControllers_21_io_II),
    .io_inConfig(configControllers_21_io_inConfig),
    .io_outConfig(configControllers_21_io_outConfig)
  );
  Dispatch_148 Dispatch_22 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_22_io_configuration),
    .io_outs_17(Dispatch_22_io_outs_17),
    .io_outs_16(Dispatch_22_io_outs_16),
    .io_outs_15(Dispatch_22_io_outs_15),
    .io_outs_14(Dispatch_22_io_outs_14),
    .io_outs_13(Dispatch_22_io_outs_13),
    .io_outs_12(Dispatch_22_io_outs_12),
    .io_outs_11(Dispatch_22_io_outs_11),
    .io_outs_10(Dispatch_22_io_outs_10),
    .io_outs_9(Dispatch_22_io_outs_9),
    .io_outs_8(Dispatch_22_io_outs_8),
    .io_outs_7(Dispatch_22_io_outs_7),
    .io_outs_6(Dispatch_22_io_outs_6),
    .io_outs_5(Dispatch_22_io_outs_5),
    .io_outs_4(Dispatch_22_io_outs_4),
    .io_outs_3(Dispatch_22_io_outs_3),
    .io_outs_2(Dispatch_22_io_outs_2),
    .io_outs_1(Dispatch_22_io_outs_1),
    .io_outs_0(Dispatch_22_io_outs_0)
  );
  ConfigController_3 configControllers_22 ( // @[TopModule.scala 262:34]
    .clock(configControllers_22_clock),
    .reset(configControllers_22_reset),
    .io_en(configControllers_22_io_en),
    .io_II(configControllers_22_io_II),
    .io_inConfig(configControllers_22_io_inConfig),
    .io_outConfig(configControllers_22_io_outConfig)
  );
  Dispatch_148 Dispatch_23 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_23_io_configuration),
    .io_outs_17(Dispatch_23_io_outs_17),
    .io_outs_16(Dispatch_23_io_outs_16),
    .io_outs_15(Dispatch_23_io_outs_15),
    .io_outs_14(Dispatch_23_io_outs_14),
    .io_outs_13(Dispatch_23_io_outs_13),
    .io_outs_12(Dispatch_23_io_outs_12),
    .io_outs_11(Dispatch_23_io_outs_11),
    .io_outs_10(Dispatch_23_io_outs_10),
    .io_outs_9(Dispatch_23_io_outs_9),
    .io_outs_8(Dispatch_23_io_outs_8),
    .io_outs_7(Dispatch_23_io_outs_7),
    .io_outs_6(Dispatch_23_io_outs_6),
    .io_outs_5(Dispatch_23_io_outs_5),
    .io_outs_4(Dispatch_23_io_outs_4),
    .io_outs_3(Dispatch_23_io_outs_3),
    .io_outs_2(Dispatch_23_io_outs_2),
    .io_outs_1(Dispatch_23_io_outs_1),
    .io_outs_0(Dispatch_23_io_outs_0)
  );
  ConfigController_3 configControllers_23 ( // @[TopModule.scala 262:34]
    .clock(configControllers_23_clock),
    .reset(configControllers_23_reset),
    .io_en(configControllers_23_io_en),
    .io_II(configControllers_23_io_II),
    .io_inConfig(configControllers_23_io_inConfig),
    .io_outConfig(configControllers_23_io_outConfig)
  );
  Dispatch_148 Dispatch_24 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_24_io_configuration),
    .io_outs_17(Dispatch_24_io_outs_17),
    .io_outs_16(Dispatch_24_io_outs_16),
    .io_outs_15(Dispatch_24_io_outs_15),
    .io_outs_14(Dispatch_24_io_outs_14),
    .io_outs_13(Dispatch_24_io_outs_13),
    .io_outs_12(Dispatch_24_io_outs_12),
    .io_outs_11(Dispatch_24_io_outs_11),
    .io_outs_10(Dispatch_24_io_outs_10),
    .io_outs_9(Dispatch_24_io_outs_9),
    .io_outs_8(Dispatch_24_io_outs_8),
    .io_outs_7(Dispatch_24_io_outs_7),
    .io_outs_6(Dispatch_24_io_outs_6),
    .io_outs_5(Dispatch_24_io_outs_5),
    .io_outs_4(Dispatch_24_io_outs_4),
    .io_outs_3(Dispatch_24_io_outs_3),
    .io_outs_2(Dispatch_24_io_outs_2),
    .io_outs_1(Dispatch_24_io_outs_1),
    .io_outs_0(Dispatch_24_io_outs_0)
  );
  ConfigController_3 configControllers_24 ( // @[TopModule.scala 262:34]
    .clock(configControllers_24_clock),
    .reset(configControllers_24_reset),
    .io_en(configControllers_24_io_en),
    .io_II(configControllers_24_io_II),
    .io_inConfig(configControllers_24_io_inConfig),
    .io_outConfig(configControllers_24_io_outConfig)
  );
  Dispatch_148 Dispatch_25 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_25_io_configuration),
    .io_outs_17(Dispatch_25_io_outs_17),
    .io_outs_16(Dispatch_25_io_outs_16),
    .io_outs_15(Dispatch_25_io_outs_15),
    .io_outs_14(Dispatch_25_io_outs_14),
    .io_outs_13(Dispatch_25_io_outs_13),
    .io_outs_12(Dispatch_25_io_outs_12),
    .io_outs_11(Dispatch_25_io_outs_11),
    .io_outs_10(Dispatch_25_io_outs_10),
    .io_outs_9(Dispatch_25_io_outs_9),
    .io_outs_8(Dispatch_25_io_outs_8),
    .io_outs_7(Dispatch_25_io_outs_7),
    .io_outs_6(Dispatch_25_io_outs_6),
    .io_outs_5(Dispatch_25_io_outs_5),
    .io_outs_4(Dispatch_25_io_outs_4),
    .io_outs_3(Dispatch_25_io_outs_3),
    .io_outs_2(Dispatch_25_io_outs_2),
    .io_outs_1(Dispatch_25_io_outs_1),
    .io_outs_0(Dispatch_25_io_outs_0)
  );
  ConfigController_2 configControllers_25 ( // @[TopModule.scala 262:34]
    .clock(configControllers_25_clock),
    .reset(configControllers_25_reset),
    .io_en(configControllers_25_io_en),
    .io_II(configControllers_25_io_II),
    .io_inConfig(configControllers_25_io_inConfig),
    .io_outConfig(configControllers_25_io_outConfig)
  );
  Dispatch_147 Dispatch_26 ( // @[TopModule.scala 267:26]
    .io_configuration(Dispatch_26_io_configuration),
    .io_outs_12(Dispatch_26_io_outs_12),
    .io_outs_11(Dispatch_26_io_outs_11),
    .io_outs_10(Dispatch_26_io_outs_10),
    .io_outs_9(Dispatch_26_io_outs_9),
    .io_outs_8(Dispatch_26_io_outs_8),
    .io_outs_7(Dispatch_26_io_outs_7),
    .io_outs_6(Dispatch_26_io_outs_6),
    .io_outs_5(Dispatch_26_io_outs_5),
    .io_outs_4(Dispatch_26_io_outs_4),
    .io_outs_3(Dispatch_26_io_outs_3),
    .io_outs_2(Dispatch_26_io_outs_2),
    .io_outs_1(Dispatch_26_io_outs_1),
    .io_outs_0(Dispatch_26_io_outs_0)
  );
  Dispatch_171 topDispatch ( // @[TopModule.scala 276:27]
    .io_configuration(topDispatch_io_configuration),
    .io_outs_25(topDispatch_io_outs_25),
    .io_outs_24(topDispatch_io_outs_24),
    .io_outs_23(topDispatch_io_outs_23),
    .io_outs_22(topDispatch_io_outs_22),
    .io_outs_21(topDispatch_io_outs_21),
    .io_outs_20(topDispatch_io_outs_20),
    .io_outs_19(topDispatch_io_outs_19),
    .io_outs_18(topDispatch_io_outs_18),
    .io_outs_17(topDispatch_io_outs_17),
    .io_outs_16(topDispatch_io_outs_16),
    .io_outs_15(topDispatch_io_outs_15),
    .io_outs_14(topDispatch_io_outs_14),
    .io_outs_13(topDispatch_io_outs_13),
    .io_outs_12(topDispatch_io_outs_12),
    .io_outs_11(topDispatch_io_outs_11),
    .io_outs_10(topDispatch_io_outs_10),
    .io_outs_9(topDispatch_io_outs_9),
    .io_outs_8(topDispatch_io_outs_8),
    .io_outs_7(topDispatch_io_outs_7),
    .io_outs_6(topDispatch_io_outs_6),
    .io_outs_5(topDispatch_io_outs_5),
    .io_outs_4(topDispatch_io_outs_4),
    .io_outs_3(topDispatch_io_outs_3),
    .io_outs_2(topDispatch_io_outs_2),
    .io_outs_1(topDispatch_io_outs_1),
    .io_outs_0(topDispatch_io_outs_0)
  );
  assign io_streamInLSU_7_ready = LoadStoreUnit_7_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_6_ready = LoadStoreUnit_6_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_5_ready = LoadStoreUnit_5_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_4_ready = LoadStoreUnit_4_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_3_ready = LoadStoreUnit_3_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_2_ready = LoadStoreUnit_2_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_1_ready = LoadStoreUnit_1_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamInLSU_0_ready = LoadStoreUnit_io_streamIn_ready; // @[TopModule.scala 195:21]
  assign io_streamOutLSU_7_valid = LoadStoreUnit_7_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_7_bits = LoadStoreUnit_7_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_6_valid = LoadStoreUnit_6_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_6_bits = LoadStoreUnit_6_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_5_valid = LoadStoreUnit_5_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_5_bits = LoadStoreUnit_5_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_4_valid = LoadStoreUnit_4_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_4_bits = LoadStoreUnit_4_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_3_valid = LoadStoreUnit_3_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_3_bits = LoadStoreUnit_3_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_2_valid = LoadStoreUnit_2_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_2_bits = LoadStoreUnit_2_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_1_valid = LoadStoreUnit_1_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_1_bits = LoadStoreUnit_1_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_0_valid = LoadStoreUnit_io_streamOut_valid; // @[TopModule.scala 196:22]
  assign io_streamOutLSU_0_bits = LoadStoreUnit_io_streamOut_bits; // @[TopModule.scala 196:22]
  assign io_idleLSU_0 = LoadStoreUnit_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_1 = LoadStoreUnit_1_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_2 = LoadStoreUnit_2_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_3 = LoadStoreUnit_3_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_4 = LoadStoreUnit_4_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_5 = LoadStoreUnit_5_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_6 = LoadStoreUnit_6_io_idle; // @[TopModule.scala 192:17]
  assign io_idleLSU_7 = LoadStoreUnit_7_io_idle; // @[TopModule.scala 192:17]
  assign io_outs_11 = RegisterFile_23_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_10 = RegisterFile_21_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_9 = RegisterFile_19_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_8 = RegisterFile_17_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_7 = RegisterFile_15_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_6 = RegisterFile_13_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_5 = RegisterFile_11_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_4 = RegisterFile_9_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_3 = RegisterFile_7_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_2 = RegisterFile_5_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_1 = RegisterFile_3_io_outs_0; // @[TopModule.scala 291:25]
  assign io_outs_0 = RegisterFile_1_io_outs_0; // @[TopModule.scala 291:25]
  assign Dispatch_io_configuration = io_schedules; // @[TopModule.scala 123:39]
  assign Alu_clock = clock;
  assign Alu_reset = reset;
  assign Alu_io_en = MultiIIScheduleController_io_valid; // @[TopModule.scala 144:17]
  assign Alu_io_skewing = MultiIIScheduleController_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_io_configuration = Dispatch_4_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_io_inputs_1 = RegisterFile_28_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_io_inputs_0 = RegisterFile_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_1_clock = clock;
  assign Alu_1_reset = reset;
  assign Alu_1_io_en = MultiIIScheduleController_1_io_valid; // @[TopModule.scala 144:17]
  assign Alu_1_io_skewing = MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_1_io_configuration = Dispatch_5_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_1_io_inputs_1 = RegisterFile_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_1_io_inputs_0 = RegisterFile_33_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_2_clock = clock;
  assign Alu_2_reset = reset;
  assign Alu_2_io_en = MultiIIScheduleController_2_io_valid; // @[TopModule.scala 144:17]
  assign Alu_2_io_skewing = MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_2_io_configuration = Dispatch_6_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_2_io_inputs_1 = RegisterFile_40_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_2_io_inputs_0 = RegisterFile_39_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_3_clock = clock;
  assign Alu_3_reset = reset;
  assign Alu_3_io_en = MultiIIScheduleController_3_io_valid; // @[TopModule.scala 144:17]
  assign Alu_3_io_skewing = MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_3_io_configuration = Dispatch_7_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_3_io_inputs_1 = RegisterFile_46_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_3_io_inputs_0 = RegisterFile_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_4_clock = clock;
  assign Alu_4_reset = reset;
  assign Alu_4_io_en = MultiIIScheduleController_4_io_valid; // @[TopModule.scala 144:17]
  assign Alu_4_io_skewing = MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_4_io_configuration = Dispatch_10_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_4_io_inputs_1 = RegisterFile_58_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_4_io_inputs_0 = RegisterFile_57_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_5_clock = clock;
  assign Alu_5_reset = reset;
  assign Alu_5_io_en = MultiIIScheduleController_5_io_valid; // @[TopModule.scala 144:17]
  assign Alu_5_io_skewing = MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_5_io_configuration = Dispatch_11_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_5_io_inputs_1 = RegisterFile_64_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_5_io_inputs_0 = RegisterFile_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_6_clock = clock;
  assign Alu_6_reset = reset;
  assign Alu_6_io_en = MultiIIScheduleController_6_io_valid; // @[TopModule.scala 144:17]
  assign Alu_6_io_skewing = MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_6_io_configuration = Dispatch_12_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_6_io_inputs_1 = RegisterFile_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_6_io_inputs_0 = RegisterFile_69_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_7_clock = clock;
  assign Alu_7_reset = reset;
  assign Alu_7_io_en = MultiIIScheduleController_7_io_valid; // @[TopModule.scala 144:17]
  assign Alu_7_io_skewing = MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_7_io_configuration = Dispatch_13_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_7_io_inputs_1 = RegisterFile_76_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_7_io_inputs_0 = RegisterFile_75_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_8_clock = clock;
  assign Alu_8_reset = reset;
  assign Alu_8_io_en = MultiIIScheduleController_8_io_valid; // @[TopModule.scala 144:17]
  assign Alu_8_io_skewing = MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_8_io_configuration = Dispatch_16_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_8_io_inputs_1 = RegisterFile_88_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_8_io_inputs_0 = RegisterFile_87_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_9_clock = clock;
  assign Alu_9_reset = reset;
  assign Alu_9_io_en = MultiIIScheduleController_9_io_valid; // @[TopModule.scala 144:17]
  assign Alu_9_io_skewing = MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_9_io_configuration = Dispatch_17_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_9_io_inputs_1 = RegisterFile_94_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_9_io_inputs_0 = RegisterFile_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_10_clock = clock;
  assign Alu_10_reset = reset;
  assign Alu_10_io_en = MultiIIScheduleController_10_io_valid; // @[TopModule.scala 144:17]
  assign Alu_10_io_skewing = MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_10_io_configuration = Dispatch_18_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_10_io_inputs_1 = RegisterFile_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_10_io_inputs_0 = RegisterFile_99_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_11_clock = clock;
  assign Alu_11_reset = reset;
  assign Alu_11_io_en = MultiIIScheduleController_11_io_valid; // @[TopModule.scala 144:17]
  assign Alu_11_io_skewing = MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_11_io_configuration = Dispatch_19_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_11_io_inputs_1 = RegisterFile_106_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_11_io_inputs_0 = RegisterFile_105_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_12_clock = clock;
  assign Alu_12_reset = reset;
  assign Alu_12_io_en = MultiIIScheduleController_12_io_valid; // @[TopModule.scala 144:17]
  assign Alu_12_io_skewing = MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_12_io_configuration = Dispatch_22_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_12_io_inputs_1 = RegisterFile_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_12_io_inputs_0 = RegisterFile_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_13_clock = clock;
  assign Alu_13_reset = reset;
  assign Alu_13_io_en = MultiIIScheduleController_13_io_valid; // @[TopModule.scala 144:17]
  assign Alu_13_io_skewing = MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_13_io_configuration = Dispatch_23_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_13_io_inputs_1 = RegisterFile_124_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_13_io_inputs_0 = RegisterFile_123_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_14_clock = clock;
  assign Alu_14_reset = reset;
  assign Alu_14_io_en = MultiIIScheduleController_14_io_valid; // @[TopModule.scala 144:17]
  assign Alu_14_io_skewing = MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_14_io_configuration = Dispatch_24_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_14_io_inputs_1 = RegisterFile_130_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_14_io_inputs_0 = RegisterFile_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_15_clock = clock;
  assign Alu_15_reset = reset;
  assign Alu_15_io_en = MultiIIScheduleController_15_io_valid; // @[TopModule.scala 144:17]
  assign Alu_15_io_skewing = MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 145:22]
  assign Alu_15_io_configuration = Dispatch_25_io_outs_0; // @[TopModule.scala 270:22]
  assign Alu_15_io_inputs_1 = RegisterFile_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Alu_15_io_inputs_0 = RegisterFile_135_io_outs_0; // @[TopModule.scala 295:60]
  assign MultiIIScheduleController_clock = clock;
  assign MultiIIScheduleController_reset = reset;
  assign MultiIIScheduleController_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_io_schedules_0 = Dispatch_io_outs_0; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_1 = Dispatch_io_outs_1; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_2 = Dispatch_io_outs_2; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_3 = Dispatch_io_outs_3; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_4 = Dispatch_io_outs_4; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_5 = Dispatch_io_outs_5; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_6 = Dispatch_io_outs_6; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_schedules_7 = Dispatch_io_outs_7; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_1_clock = clock;
  assign MultiIIScheduleController_1_reset = reset;
  assign MultiIIScheduleController_1_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_1_io_schedules_0 = Dispatch_io_outs_8; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_1 = Dispatch_io_outs_9; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_2 = Dispatch_io_outs_10; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_3 = Dispatch_io_outs_11; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_4 = Dispatch_io_outs_12; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_5 = Dispatch_io_outs_13; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_6 = Dispatch_io_outs_14; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_schedules_7 = Dispatch_io_outs_15; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_1_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_2_clock = clock;
  assign MultiIIScheduleController_2_reset = reset;
  assign MultiIIScheduleController_2_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_2_io_schedules_0 = Dispatch_io_outs_16; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_1 = Dispatch_io_outs_17; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_2 = Dispatch_io_outs_18; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_3 = Dispatch_io_outs_19; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_4 = Dispatch_io_outs_20; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_5 = Dispatch_io_outs_21; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_6 = Dispatch_io_outs_22; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_schedules_7 = Dispatch_io_outs_23; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_2_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_3_clock = clock;
  assign MultiIIScheduleController_3_reset = reset;
  assign MultiIIScheduleController_3_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_3_io_schedules_0 = Dispatch_io_outs_24; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_1 = Dispatch_io_outs_25; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_2 = Dispatch_io_outs_26; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_3 = Dispatch_io_outs_27; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_4 = Dispatch_io_outs_28; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_5 = Dispatch_io_outs_29; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_6 = Dispatch_io_outs_30; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_schedules_7 = Dispatch_io_outs_31; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_3_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_4_clock = clock;
  assign MultiIIScheduleController_4_reset = reset;
  assign MultiIIScheduleController_4_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_4_io_schedules_0 = Dispatch_io_outs_32; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_1 = Dispatch_io_outs_33; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_2 = Dispatch_io_outs_34; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_3 = Dispatch_io_outs_35; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_4 = Dispatch_io_outs_36; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_5 = Dispatch_io_outs_37; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_6 = Dispatch_io_outs_38; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_schedules_7 = Dispatch_io_outs_39; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_4_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_5_clock = clock;
  assign MultiIIScheduleController_5_reset = reset;
  assign MultiIIScheduleController_5_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_5_io_schedules_0 = Dispatch_io_outs_40; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_1 = Dispatch_io_outs_41; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_2 = Dispatch_io_outs_42; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_3 = Dispatch_io_outs_43; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_4 = Dispatch_io_outs_44; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_5 = Dispatch_io_outs_45; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_6 = Dispatch_io_outs_46; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_schedules_7 = Dispatch_io_outs_47; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_5_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_6_clock = clock;
  assign MultiIIScheduleController_6_reset = reset;
  assign MultiIIScheduleController_6_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_6_io_schedules_0 = Dispatch_io_outs_48; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_1 = Dispatch_io_outs_49; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_2 = Dispatch_io_outs_50; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_3 = Dispatch_io_outs_51; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_4 = Dispatch_io_outs_52; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_5 = Dispatch_io_outs_53; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_6 = Dispatch_io_outs_54; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_schedules_7 = Dispatch_io_outs_55; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_6_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_7_clock = clock;
  assign MultiIIScheduleController_7_reset = reset;
  assign MultiIIScheduleController_7_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_7_io_schedules_0 = Dispatch_io_outs_56; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_1 = Dispatch_io_outs_57; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_2 = Dispatch_io_outs_58; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_3 = Dispatch_io_outs_59; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_4 = Dispatch_io_outs_60; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_5 = Dispatch_io_outs_61; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_6 = Dispatch_io_outs_62; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_schedules_7 = Dispatch_io_outs_63; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_7_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_8_clock = clock;
  assign MultiIIScheduleController_8_reset = reset;
  assign MultiIIScheduleController_8_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_8_io_schedules_0 = Dispatch_io_outs_64; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_1 = Dispatch_io_outs_65; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_2 = Dispatch_io_outs_66; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_3 = Dispatch_io_outs_67; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_4 = Dispatch_io_outs_68; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_5 = Dispatch_io_outs_69; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_6 = Dispatch_io_outs_70; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_schedules_7 = Dispatch_io_outs_71; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_8_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_9_clock = clock;
  assign MultiIIScheduleController_9_reset = reset;
  assign MultiIIScheduleController_9_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_9_io_schedules_0 = Dispatch_io_outs_72; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_1 = Dispatch_io_outs_73; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_2 = Dispatch_io_outs_74; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_3 = Dispatch_io_outs_75; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_4 = Dispatch_io_outs_76; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_5 = Dispatch_io_outs_77; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_6 = Dispatch_io_outs_78; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_schedules_7 = Dispatch_io_outs_79; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_9_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_10_clock = clock;
  assign MultiIIScheduleController_10_reset = reset;
  assign MultiIIScheduleController_10_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_10_io_schedules_0 = Dispatch_io_outs_80; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_1 = Dispatch_io_outs_81; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_2 = Dispatch_io_outs_82; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_3 = Dispatch_io_outs_83; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_4 = Dispatch_io_outs_84; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_5 = Dispatch_io_outs_85; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_6 = Dispatch_io_outs_86; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_schedules_7 = Dispatch_io_outs_87; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_10_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_11_clock = clock;
  assign MultiIIScheduleController_11_reset = reset;
  assign MultiIIScheduleController_11_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_11_io_schedules_0 = Dispatch_io_outs_88; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_1 = Dispatch_io_outs_89; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_2 = Dispatch_io_outs_90; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_3 = Dispatch_io_outs_91; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_4 = Dispatch_io_outs_92; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_5 = Dispatch_io_outs_93; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_6 = Dispatch_io_outs_94; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_schedules_7 = Dispatch_io_outs_95; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_11_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_12_clock = clock;
  assign MultiIIScheduleController_12_reset = reset;
  assign MultiIIScheduleController_12_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_12_io_schedules_0 = Dispatch_io_outs_96; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_1 = Dispatch_io_outs_97; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_2 = Dispatch_io_outs_98; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_3 = Dispatch_io_outs_99; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_4 = Dispatch_io_outs_100; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_5 = Dispatch_io_outs_101; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_6 = Dispatch_io_outs_102; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_schedules_7 = Dispatch_io_outs_103; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_12_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_13_clock = clock;
  assign MultiIIScheduleController_13_reset = reset;
  assign MultiIIScheduleController_13_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_13_io_schedules_0 = Dispatch_io_outs_104; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_1 = Dispatch_io_outs_105; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_2 = Dispatch_io_outs_106; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_3 = Dispatch_io_outs_107; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_4 = Dispatch_io_outs_108; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_5 = Dispatch_io_outs_109; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_6 = Dispatch_io_outs_110; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_schedules_7 = Dispatch_io_outs_111; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_13_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_14_clock = clock;
  assign MultiIIScheduleController_14_reset = reset;
  assign MultiIIScheduleController_14_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_14_io_schedules_0 = Dispatch_io_outs_112; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_1 = Dispatch_io_outs_113; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_2 = Dispatch_io_outs_114; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_3 = Dispatch_io_outs_115; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_4 = Dispatch_io_outs_116; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_5 = Dispatch_io_outs_117; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_6 = Dispatch_io_outs_118; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_schedules_7 = Dispatch_io_outs_119; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_14_io_II = io_II; // @[TopModule.scala 140:35]
  assign MultiIIScheduleController_15_clock = clock;
  assign MultiIIScheduleController_15_reset = reset;
  assign MultiIIScheduleController_15_io_en = io_en; // @[TopModule.scala 139:35]
  assign MultiIIScheduleController_15_io_schedules_0 = Dispatch_io_outs_120; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_1 = Dispatch_io_outs_121; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_2 = Dispatch_io_outs_122; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_3 = Dispatch_io_outs_123; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_4 = Dispatch_io_outs_124; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_5 = Dispatch_io_outs_125; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_6 = Dispatch_io_outs_126; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_schedules_7 = Dispatch_io_outs_127; // @[TopModule.scala 142:47]
  assign MultiIIScheduleController_15_io_II = io_II; // @[TopModule.scala 140:35]
  assign RegisterFile_clock = clock;
  assign RegisterFile_reset = reset;
  assign RegisterFile_io_configuration = Dispatch_1_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_io_inputs_0 = io_inputs_0; // @[TopModule.scala 293:60]
  assign RegisterFile_1_clock = clock;
  assign RegisterFile_1_reset = reset;
  assign RegisterFile_1_io_configuration = Dispatch_1_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_1_io_inputs_0 = Multiplexer_6_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_2_clock = clock;
  assign RegisterFile_2_reset = reset;
  assign RegisterFile_2_io_configuration = Dispatch_1_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_2_io_inputs_0 = io_inputs_1; // @[TopModule.scala 293:60]
  assign RegisterFile_3_clock = clock;
  assign RegisterFile_3_reset = reset;
  assign RegisterFile_3_io_configuration = Dispatch_1_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_3_io_inputs_0 = Multiplexer_16_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_4_clock = clock;
  assign RegisterFile_4_reset = reset;
  assign RegisterFile_4_io_configuration = Dispatch_1_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_4_io_inputs_0 = io_inputs_2; // @[TopModule.scala 293:60]
  assign RegisterFile_5_clock = clock;
  assign RegisterFile_5_reset = reset;
  assign RegisterFile_5_io_configuration = Dispatch_1_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_5_io_inputs_0 = Multiplexer_26_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_6_clock = clock;
  assign RegisterFile_6_reset = reset;
  assign RegisterFile_6_io_configuration = Dispatch_1_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_6_io_inputs_0 = io_inputs_3; // @[TopModule.scala 293:60]
  assign RegisterFile_7_clock = clock;
  assign RegisterFile_7_reset = reset;
  assign RegisterFile_7_io_configuration = Dispatch_1_io_outs_7; // @[TopModule.scala 270:22]
  assign RegisterFile_7_io_inputs_0 = Multiplexer_36_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_8_clock = clock;
  assign RegisterFile_8_reset = reset;
  assign RegisterFile_8_io_configuration = Dispatch_1_io_outs_8; // @[TopModule.scala 270:22]
  assign RegisterFile_8_io_inputs_0 = io_inputs_4; // @[TopModule.scala 293:60]
  assign RegisterFile_9_clock = clock;
  assign RegisterFile_9_reset = reset;
  assign RegisterFile_9_io_configuration = Dispatch_1_io_outs_9; // @[TopModule.scala 270:22]
  assign RegisterFile_9_io_inputs_0 = Multiplexer_46_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_10_clock = clock;
  assign RegisterFile_10_reset = reset;
  assign RegisterFile_10_io_configuration = Dispatch_1_io_outs_10; // @[TopModule.scala 270:22]
  assign RegisterFile_10_io_inputs_0 = io_inputs_5; // @[TopModule.scala 293:60]
  assign RegisterFile_11_clock = clock;
  assign RegisterFile_11_reset = reset;
  assign RegisterFile_11_io_configuration = Dispatch_1_io_outs_11; // @[TopModule.scala 270:22]
  assign RegisterFile_11_io_inputs_0 = Multiplexer_55_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_12_clock = clock;
  assign RegisterFile_12_reset = reset;
  assign RegisterFile_12_io_configuration = Dispatch_2_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_12_io_inputs_0 = io_inputs_6; // @[TopModule.scala 293:60]
  assign RegisterFile_13_clock = clock;
  assign RegisterFile_13_reset = reset;
  assign RegisterFile_13_io_configuration = Dispatch_2_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_13_io_inputs_0 = Multiplexer_174_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_14_clock = clock;
  assign RegisterFile_14_reset = reset;
  assign RegisterFile_14_io_configuration = Dispatch_2_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_14_io_inputs_0 = io_inputs_7; // @[TopModule.scala 293:60]
  assign RegisterFile_15_clock = clock;
  assign RegisterFile_15_reset = reset;
  assign RegisterFile_15_io_configuration = Dispatch_2_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_15_io_inputs_0 = Multiplexer_184_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_16_clock = clock;
  assign RegisterFile_16_reset = reset;
  assign RegisterFile_16_io_configuration = Dispatch_2_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_16_io_inputs_0 = io_inputs_8; // @[TopModule.scala 293:60]
  assign RegisterFile_17_clock = clock;
  assign RegisterFile_17_reset = reset;
  assign RegisterFile_17_io_configuration = Dispatch_2_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_17_io_inputs_0 = Multiplexer_194_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_18_clock = clock;
  assign RegisterFile_18_reset = reset;
  assign RegisterFile_18_io_configuration = Dispatch_2_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_18_io_inputs_0 = io_inputs_9; // @[TopModule.scala 293:60]
  assign RegisterFile_19_clock = clock;
  assign RegisterFile_19_reset = reset;
  assign RegisterFile_19_io_configuration = Dispatch_2_io_outs_7; // @[TopModule.scala 270:22]
  assign RegisterFile_19_io_inputs_0 = Multiplexer_204_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_20_clock = clock;
  assign RegisterFile_20_reset = reset;
  assign RegisterFile_20_io_configuration = Dispatch_2_io_outs_8; // @[TopModule.scala 270:22]
  assign RegisterFile_20_io_inputs_0 = io_inputs_10; // @[TopModule.scala 293:60]
  assign RegisterFile_21_clock = clock;
  assign RegisterFile_21_reset = reset;
  assign RegisterFile_21_io_configuration = Dispatch_2_io_outs_9; // @[TopModule.scala 270:22]
  assign RegisterFile_21_io_inputs_0 = Multiplexer_214_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_22_clock = clock;
  assign RegisterFile_22_reset = reset;
  assign RegisterFile_22_io_configuration = Dispatch_2_io_outs_10; // @[TopModule.scala 270:22]
  assign RegisterFile_22_io_inputs_0 = io_inputs_11; // @[TopModule.scala 293:60]
  assign RegisterFile_23_clock = clock;
  assign RegisterFile_23_reset = reset;
  assign RegisterFile_23_io_configuration = Dispatch_2_io_outs_11; // @[TopModule.scala 270:22]
  assign RegisterFile_23_io_inputs_0 = Multiplexer_223_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_24_clock = clock;
  assign RegisterFile_24_reset = reset;
  assign RegisterFile_24_io_configuration = Dispatch_3_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_24_io_inputs_0 = Multiplexer_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_25_clock = clock;
  assign RegisterFile_25_reset = reset;
  assign RegisterFile_25_io_configuration = Dispatch_3_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_25_io_inputs_0 = Multiplexer_1_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_26_clock = clock;
  assign RegisterFile_26_reset = reset;
  assign RegisterFile_26_io_configuration = Dispatch_3_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_26_io_inputs_0 = Multiplexer_2_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_27_clock = clock;
  assign RegisterFile_27_reset = reset;
  assign RegisterFile_27_io_configuration = Dispatch_4_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_27_io_inputs_0 = Multiplexer_12_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_28_clock = clock;
  assign RegisterFile_28_reset = reset;
  assign RegisterFile_28_io_configuration = Dispatch_4_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_28_io_inputs_0 = Multiplexer_13_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_29_clock = clock;
  assign RegisterFile_29_reset = reset;
  assign RegisterFile_29_io_configuration = Dispatch_4_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_29_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_30_clock = clock;
  assign RegisterFile_30_reset = reset;
  assign RegisterFile_30_io_configuration = Dispatch_4_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_30_io_inputs_0 = Multiplexer_9_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_31_clock = clock;
  assign RegisterFile_31_reset = reset;
  assign RegisterFile_31_io_configuration = Dispatch_4_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_31_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_32_clock = clock;
  assign RegisterFile_32_reset = reset;
  assign RegisterFile_32_io_configuration = Dispatch_4_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_32_io_inputs_0 = Multiplexer_11_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_33_clock = clock;
  assign RegisterFile_33_reset = reset;
  assign RegisterFile_33_io_configuration = Dispatch_5_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_33_io_inputs_0 = Multiplexer_22_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_34_clock = clock;
  assign RegisterFile_34_reset = reset;
  assign RegisterFile_34_io_configuration = Dispatch_5_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_34_io_inputs_0 = Multiplexer_23_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_35_clock = clock;
  assign RegisterFile_35_reset = reset;
  assign RegisterFile_35_io_configuration = Dispatch_5_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_35_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_36_clock = clock;
  assign RegisterFile_36_reset = reset;
  assign RegisterFile_36_io_configuration = Dispatch_5_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_36_io_inputs_0 = Multiplexer_19_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_37_clock = clock;
  assign RegisterFile_37_reset = reset;
  assign RegisterFile_37_io_configuration = Dispatch_5_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_37_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_38_clock = clock;
  assign RegisterFile_38_reset = reset;
  assign RegisterFile_38_io_configuration = Dispatch_5_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_38_io_inputs_0 = Multiplexer_21_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_39_clock = clock;
  assign RegisterFile_39_reset = reset;
  assign RegisterFile_39_io_configuration = Dispatch_6_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_39_io_inputs_0 = Multiplexer_32_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_40_clock = clock;
  assign RegisterFile_40_reset = reset;
  assign RegisterFile_40_io_configuration = Dispatch_6_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_40_io_inputs_0 = Multiplexer_33_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_41_clock = clock;
  assign RegisterFile_41_reset = reset;
  assign RegisterFile_41_io_configuration = Dispatch_6_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_41_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_42_clock = clock;
  assign RegisterFile_42_reset = reset;
  assign RegisterFile_42_io_configuration = Dispatch_6_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_42_io_inputs_0 = Multiplexer_29_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_43_clock = clock;
  assign RegisterFile_43_reset = reset;
  assign RegisterFile_43_io_configuration = Dispatch_6_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_43_io_inputs_0 = Multiplexer_30_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_44_clock = clock;
  assign RegisterFile_44_reset = reset;
  assign RegisterFile_44_io_configuration = Dispatch_6_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_44_io_inputs_0 = Multiplexer_31_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_45_clock = clock;
  assign RegisterFile_45_reset = reset;
  assign RegisterFile_45_io_configuration = Dispatch_7_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_45_io_inputs_0 = Multiplexer_42_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_46_clock = clock;
  assign RegisterFile_46_reset = reset;
  assign RegisterFile_46_io_configuration = Dispatch_7_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_46_io_inputs_0 = Multiplexer_43_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_47_clock = clock;
  assign RegisterFile_47_reset = reset;
  assign RegisterFile_47_io_configuration = Dispatch_7_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_47_io_inputs_0 = Multiplexer_38_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_48_clock = clock;
  assign RegisterFile_48_reset = reset;
  assign RegisterFile_48_io_configuration = Dispatch_7_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_48_io_inputs_0 = Multiplexer_39_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_49_clock = clock;
  assign RegisterFile_49_reset = reset;
  assign RegisterFile_49_io_configuration = Dispatch_7_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_49_io_inputs_0 = Multiplexer_40_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_50_clock = clock;
  assign RegisterFile_50_reset = reset;
  assign RegisterFile_50_io_configuration = Dispatch_7_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_50_io_inputs_0 = Multiplexer_41_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_51_clock = clock;
  assign RegisterFile_51_reset = reset;
  assign RegisterFile_51_io_configuration = Dispatch_8_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_51_io_inputs_0 = Multiplexer_48_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_52_clock = clock;
  assign RegisterFile_52_reset = reset;
  assign RegisterFile_52_io_configuration = Dispatch_8_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_52_io_inputs_0 = Multiplexer_49_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_53_clock = clock;
  assign RegisterFile_53_reset = reset;
  assign RegisterFile_53_io_configuration = Dispatch_8_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_53_io_inputs_0 = Multiplexer_50_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_54_clock = clock;
  assign RegisterFile_54_reset = reset;
  assign RegisterFile_54_io_configuration = Dispatch_9_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_54_io_inputs_0 = Multiplexer_56_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_55_clock = clock;
  assign RegisterFile_55_reset = reset;
  assign RegisterFile_55_io_configuration = Dispatch_9_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_55_io_inputs_0 = Multiplexer_57_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_56_clock = clock;
  assign RegisterFile_56_reset = reset;
  assign RegisterFile_56_io_configuration = Dispatch_9_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_56_io_inputs_0 = Multiplexer_58_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_57_clock = clock;
  assign RegisterFile_57_reset = reset;
  assign RegisterFile_57_io_configuration = Dispatch_10_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_57_io_inputs_0 = Multiplexer_68_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_58_clock = clock;
  assign RegisterFile_58_reset = reset;
  assign RegisterFile_58_io_configuration = Dispatch_10_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_58_io_inputs_0 = Multiplexer_69_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_59_clock = clock;
  assign RegisterFile_59_reset = reset;
  assign RegisterFile_59_io_configuration = Dispatch_10_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_59_io_inputs_0 = Multiplexer_64_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_60_clock = clock;
  assign RegisterFile_60_reset = reset;
  assign RegisterFile_60_io_configuration = Dispatch_10_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_60_io_inputs_0 = Multiplexer_65_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_61_clock = clock;
  assign RegisterFile_61_reset = reset;
  assign RegisterFile_61_io_configuration = Dispatch_10_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_61_io_inputs_0 = Multiplexer_66_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_62_clock = clock;
  assign RegisterFile_62_reset = reset;
  assign RegisterFile_62_io_configuration = Dispatch_10_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_62_io_inputs_0 = Multiplexer_67_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_63_clock = clock;
  assign RegisterFile_63_reset = reset;
  assign RegisterFile_63_io_configuration = Dispatch_11_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_63_io_inputs_0 = Multiplexer_78_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_64_clock = clock;
  assign RegisterFile_64_reset = reset;
  assign RegisterFile_64_io_configuration = Dispatch_11_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_64_io_inputs_0 = Multiplexer_79_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_65_clock = clock;
  assign RegisterFile_65_reset = reset;
  assign RegisterFile_65_io_configuration = Dispatch_11_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_65_io_inputs_0 = Multiplexer_74_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_66_clock = clock;
  assign RegisterFile_66_reset = reset;
  assign RegisterFile_66_io_configuration = Dispatch_11_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_66_io_inputs_0 = Multiplexer_75_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_67_clock = clock;
  assign RegisterFile_67_reset = reset;
  assign RegisterFile_67_io_configuration = Dispatch_11_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_67_io_inputs_0 = Multiplexer_76_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_68_clock = clock;
  assign RegisterFile_68_reset = reset;
  assign RegisterFile_68_io_configuration = Dispatch_11_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_68_io_inputs_0 = Multiplexer_77_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_69_clock = clock;
  assign RegisterFile_69_reset = reset;
  assign RegisterFile_69_io_configuration = Dispatch_12_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_69_io_inputs_0 = Multiplexer_88_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_70_clock = clock;
  assign RegisterFile_70_reset = reset;
  assign RegisterFile_70_io_configuration = Dispatch_12_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_70_io_inputs_0 = Multiplexer_89_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_71_clock = clock;
  assign RegisterFile_71_reset = reset;
  assign RegisterFile_71_io_configuration = Dispatch_12_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_71_io_inputs_0 = Multiplexer_84_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_72_clock = clock;
  assign RegisterFile_72_reset = reset;
  assign RegisterFile_72_io_configuration = Dispatch_12_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_72_io_inputs_0 = Multiplexer_85_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_73_clock = clock;
  assign RegisterFile_73_reset = reset;
  assign RegisterFile_73_io_configuration = Dispatch_12_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_73_io_inputs_0 = Multiplexer_86_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_74_clock = clock;
  assign RegisterFile_74_reset = reset;
  assign RegisterFile_74_io_configuration = Dispatch_12_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_74_io_inputs_0 = Multiplexer_87_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_75_clock = clock;
  assign RegisterFile_75_reset = reset;
  assign RegisterFile_75_io_configuration = Dispatch_13_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_75_io_inputs_0 = Multiplexer_98_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_76_clock = clock;
  assign RegisterFile_76_reset = reset;
  assign RegisterFile_76_io_configuration = Dispatch_13_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_76_io_inputs_0 = Multiplexer_99_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_77_clock = clock;
  assign RegisterFile_77_reset = reset;
  assign RegisterFile_77_io_configuration = Dispatch_13_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_77_io_inputs_0 = Multiplexer_94_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_78_clock = clock;
  assign RegisterFile_78_reset = reset;
  assign RegisterFile_78_io_configuration = Dispatch_13_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_78_io_inputs_0 = Multiplexer_95_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_79_clock = clock;
  assign RegisterFile_79_reset = reset;
  assign RegisterFile_79_io_configuration = Dispatch_13_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_79_io_inputs_0 = Multiplexer_96_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_80_clock = clock;
  assign RegisterFile_80_reset = reset;
  assign RegisterFile_80_io_configuration = Dispatch_13_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_80_io_inputs_0 = Multiplexer_97_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_81_clock = clock;
  assign RegisterFile_81_reset = reset;
  assign RegisterFile_81_io_configuration = Dispatch_14_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_81_io_inputs_0 = Multiplexer_104_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_82_clock = clock;
  assign RegisterFile_82_reset = reset;
  assign RegisterFile_82_io_configuration = Dispatch_14_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_82_io_inputs_0 = Multiplexer_105_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_83_clock = clock;
  assign RegisterFile_83_reset = reset;
  assign RegisterFile_83_io_configuration = Dispatch_14_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_83_io_inputs_0 = Multiplexer_106_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_84_clock = clock;
  assign RegisterFile_84_reset = reset;
  assign RegisterFile_84_io_configuration = Dispatch_15_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_84_io_inputs_0 = Multiplexer_112_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_85_clock = clock;
  assign RegisterFile_85_reset = reset;
  assign RegisterFile_85_io_configuration = Dispatch_15_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_85_io_inputs_0 = Multiplexer_113_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_86_clock = clock;
  assign RegisterFile_86_reset = reset;
  assign RegisterFile_86_io_configuration = Dispatch_15_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_86_io_inputs_0 = Multiplexer_114_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_87_clock = clock;
  assign RegisterFile_87_reset = reset;
  assign RegisterFile_87_io_configuration = Dispatch_16_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_87_io_inputs_0 = Multiplexer_124_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_88_clock = clock;
  assign RegisterFile_88_reset = reset;
  assign RegisterFile_88_io_configuration = Dispatch_16_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_88_io_inputs_0 = Multiplexer_125_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_89_clock = clock;
  assign RegisterFile_89_reset = reset;
  assign RegisterFile_89_io_configuration = Dispatch_16_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_89_io_inputs_0 = Multiplexer_120_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_90_clock = clock;
  assign RegisterFile_90_reset = reset;
  assign RegisterFile_90_io_configuration = Dispatch_16_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_90_io_inputs_0 = Multiplexer_121_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_91_clock = clock;
  assign RegisterFile_91_reset = reset;
  assign RegisterFile_91_io_configuration = Dispatch_16_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_91_io_inputs_0 = Multiplexer_122_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_92_clock = clock;
  assign RegisterFile_92_reset = reset;
  assign RegisterFile_92_io_configuration = Dispatch_16_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_92_io_inputs_0 = Multiplexer_123_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_93_clock = clock;
  assign RegisterFile_93_reset = reset;
  assign RegisterFile_93_io_configuration = Dispatch_17_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_93_io_inputs_0 = Multiplexer_134_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_94_clock = clock;
  assign RegisterFile_94_reset = reset;
  assign RegisterFile_94_io_configuration = Dispatch_17_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_94_io_inputs_0 = Multiplexer_135_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_95_clock = clock;
  assign RegisterFile_95_reset = reset;
  assign RegisterFile_95_io_configuration = Dispatch_17_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_95_io_inputs_0 = Multiplexer_130_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_96_clock = clock;
  assign RegisterFile_96_reset = reset;
  assign RegisterFile_96_io_configuration = Dispatch_17_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_96_io_inputs_0 = Multiplexer_131_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_97_clock = clock;
  assign RegisterFile_97_reset = reset;
  assign RegisterFile_97_io_configuration = Dispatch_17_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_97_io_inputs_0 = Multiplexer_132_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_98_clock = clock;
  assign RegisterFile_98_reset = reset;
  assign RegisterFile_98_io_configuration = Dispatch_17_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_98_io_inputs_0 = Multiplexer_133_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_99_clock = clock;
  assign RegisterFile_99_reset = reset;
  assign RegisterFile_99_io_configuration = Dispatch_18_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_99_io_inputs_0 = Multiplexer_144_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_100_clock = clock;
  assign RegisterFile_100_reset = reset;
  assign RegisterFile_100_io_configuration = Dispatch_18_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_100_io_inputs_0 = Multiplexer_145_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_101_clock = clock;
  assign RegisterFile_101_reset = reset;
  assign RegisterFile_101_io_configuration = Dispatch_18_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_101_io_inputs_0 = Multiplexer_140_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_102_clock = clock;
  assign RegisterFile_102_reset = reset;
  assign RegisterFile_102_io_configuration = Dispatch_18_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_102_io_inputs_0 = Multiplexer_141_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_103_clock = clock;
  assign RegisterFile_103_reset = reset;
  assign RegisterFile_103_io_configuration = Dispatch_18_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_103_io_inputs_0 = Multiplexer_142_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_104_clock = clock;
  assign RegisterFile_104_reset = reset;
  assign RegisterFile_104_io_configuration = Dispatch_18_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_104_io_inputs_0 = Multiplexer_143_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_105_clock = clock;
  assign RegisterFile_105_reset = reset;
  assign RegisterFile_105_io_configuration = Dispatch_19_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_105_io_inputs_0 = Multiplexer_154_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_106_clock = clock;
  assign RegisterFile_106_reset = reset;
  assign RegisterFile_106_io_configuration = Dispatch_19_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_106_io_inputs_0 = Multiplexer_155_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_107_clock = clock;
  assign RegisterFile_107_reset = reset;
  assign RegisterFile_107_io_configuration = Dispatch_19_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_107_io_inputs_0 = Multiplexer_150_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_108_clock = clock;
  assign RegisterFile_108_reset = reset;
  assign RegisterFile_108_io_configuration = Dispatch_19_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_108_io_inputs_0 = Multiplexer_151_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_109_clock = clock;
  assign RegisterFile_109_reset = reset;
  assign RegisterFile_109_io_configuration = Dispatch_19_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_109_io_inputs_0 = Multiplexer_152_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_110_clock = clock;
  assign RegisterFile_110_reset = reset;
  assign RegisterFile_110_io_configuration = Dispatch_19_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_110_io_inputs_0 = Multiplexer_153_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_111_clock = clock;
  assign RegisterFile_111_reset = reset;
  assign RegisterFile_111_io_configuration = Dispatch_20_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_111_io_inputs_0 = Multiplexer_160_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_112_clock = clock;
  assign RegisterFile_112_reset = reset;
  assign RegisterFile_112_io_configuration = Dispatch_20_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_112_io_inputs_0 = Multiplexer_161_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_113_clock = clock;
  assign RegisterFile_113_reset = reset;
  assign RegisterFile_113_io_configuration = Dispatch_20_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_113_io_inputs_0 = Multiplexer_162_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_114_clock = clock;
  assign RegisterFile_114_reset = reset;
  assign RegisterFile_114_io_configuration = Dispatch_21_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_114_io_inputs_0 = Multiplexer_168_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_115_clock = clock;
  assign RegisterFile_115_reset = reset;
  assign RegisterFile_115_io_configuration = Dispatch_21_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_115_io_inputs_0 = Multiplexer_169_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_116_clock = clock;
  assign RegisterFile_116_reset = reset;
  assign RegisterFile_116_io_configuration = Dispatch_21_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_116_io_inputs_0 = Multiplexer_170_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_117_clock = clock;
  assign RegisterFile_117_reset = reset;
  assign RegisterFile_117_io_configuration = Dispatch_22_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_117_io_inputs_0 = Multiplexer_180_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_118_clock = clock;
  assign RegisterFile_118_reset = reset;
  assign RegisterFile_118_io_configuration = Dispatch_22_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_118_io_inputs_0 = Multiplexer_181_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_119_clock = clock;
  assign RegisterFile_119_reset = reset;
  assign RegisterFile_119_io_configuration = Dispatch_22_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_119_io_inputs_0 = Multiplexer_176_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_120_clock = clock;
  assign RegisterFile_120_reset = reset;
  assign RegisterFile_120_io_configuration = Dispatch_22_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_120_io_inputs_0 = Multiplexer_177_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_121_clock = clock;
  assign RegisterFile_121_reset = reset;
  assign RegisterFile_121_io_configuration = Dispatch_22_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_121_io_inputs_0 = Multiplexer_178_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_122_clock = clock;
  assign RegisterFile_122_reset = reset;
  assign RegisterFile_122_io_configuration = Dispatch_22_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_122_io_inputs_0 = Multiplexer_179_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_123_clock = clock;
  assign RegisterFile_123_reset = reset;
  assign RegisterFile_123_io_configuration = Dispatch_23_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_123_io_inputs_0 = Multiplexer_190_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_124_clock = clock;
  assign RegisterFile_124_reset = reset;
  assign RegisterFile_124_io_configuration = Dispatch_23_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_124_io_inputs_0 = Multiplexer_191_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_125_clock = clock;
  assign RegisterFile_125_reset = reset;
  assign RegisterFile_125_io_configuration = Dispatch_23_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_125_io_inputs_0 = Multiplexer_186_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_126_clock = clock;
  assign RegisterFile_126_reset = reset;
  assign RegisterFile_126_io_configuration = Dispatch_23_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_126_io_inputs_0 = Multiplexer_187_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_127_clock = clock;
  assign RegisterFile_127_reset = reset;
  assign RegisterFile_127_io_configuration = Dispatch_23_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_127_io_inputs_0 = Multiplexer_188_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_128_clock = clock;
  assign RegisterFile_128_reset = reset;
  assign RegisterFile_128_io_configuration = Dispatch_23_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_128_io_inputs_0 = Multiplexer_189_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_129_clock = clock;
  assign RegisterFile_129_reset = reset;
  assign RegisterFile_129_io_configuration = Dispatch_24_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_129_io_inputs_0 = Multiplexer_200_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_130_clock = clock;
  assign RegisterFile_130_reset = reset;
  assign RegisterFile_130_io_configuration = Dispatch_24_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_130_io_inputs_0 = Multiplexer_201_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_131_clock = clock;
  assign RegisterFile_131_reset = reset;
  assign RegisterFile_131_io_configuration = Dispatch_24_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_131_io_inputs_0 = Multiplexer_196_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_132_clock = clock;
  assign RegisterFile_132_reset = reset;
  assign RegisterFile_132_io_configuration = Dispatch_24_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_132_io_inputs_0 = Multiplexer_197_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_133_clock = clock;
  assign RegisterFile_133_reset = reset;
  assign RegisterFile_133_io_configuration = Dispatch_24_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_133_io_inputs_0 = Multiplexer_198_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_134_clock = clock;
  assign RegisterFile_134_reset = reset;
  assign RegisterFile_134_io_configuration = Dispatch_24_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_134_io_inputs_0 = Multiplexer_199_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_135_clock = clock;
  assign RegisterFile_135_reset = reset;
  assign RegisterFile_135_io_configuration = Dispatch_25_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_135_io_inputs_0 = Multiplexer_210_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_136_clock = clock;
  assign RegisterFile_136_reset = reset;
  assign RegisterFile_136_io_configuration = Dispatch_25_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_136_io_inputs_0 = Multiplexer_211_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_137_clock = clock;
  assign RegisterFile_137_reset = reset;
  assign RegisterFile_137_io_configuration = Dispatch_25_io_outs_3; // @[TopModule.scala 270:22]
  assign RegisterFile_137_io_inputs_0 = Multiplexer_206_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_138_clock = clock;
  assign RegisterFile_138_reset = reset;
  assign RegisterFile_138_io_configuration = Dispatch_25_io_outs_4; // @[TopModule.scala 270:22]
  assign RegisterFile_138_io_inputs_0 = Multiplexer_207_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_139_clock = clock;
  assign RegisterFile_139_reset = reset;
  assign RegisterFile_139_io_configuration = Dispatch_25_io_outs_5; // @[TopModule.scala 270:22]
  assign RegisterFile_139_io_inputs_0 = Multiplexer_208_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_140_clock = clock;
  assign RegisterFile_140_reset = reset;
  assign RegisterFile_140_io_configuration = Dispatch_25_io_outs_6; // @[TopModule.scala 270:22]
  assign RegisterFile_140_io_inputs_0 = Multiplexer_209_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_141_clock = clock;
  assign RegisterFile_141_reset = reset;
  assign RegisterFile_141_io_configuration = Dispatch_26_io_outs_0; // @[TopModule.scala 270:22]
  assign RegisterFile_141_io_inputs_0 = Multiplexer_216_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_142_clock = clock;
  assign RegisterFile_142_reset = reset;
  assign RegisterFile_142_io_configuration = Dispatch_26_io_outs_1; // @[TopModule.scala 270:22]
  assign RegisterFile_142_io_inputs_0 = Multiplexer_217_io_outs_0; // @[TopModule.scala 295:60]
  assign RegisterFile_143_clock = clock;
  assign RegisterFile_143_reset = reset;
  assign RegisterFile_143_io_configuration = Dispatch_26_io_outs_2; // @[TopModule.scala 270:22]
  assign RegisterFile_143_io_inputs_0 = Multiplexer_218_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_io_configuration = Dispatch_3_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_io_inputs_3 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_io_inputs_2 = Multiplexer_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_io_inputs_1 = RegisterFile_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_io_inputs_0 = Multiplexer_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_1_io_configuration = Dispatch_3_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_1_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_1_io_inputs_3 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_1_io_inputs_2 = Multiplexer_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_1_io_inputs_1 = RegisterFile_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_1_io_inputs_0 = Multiplexer_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_2_io_configuration = Dispatch_3_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_2_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_2_io_inputs_3 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_2_io_inputs_2 = Multiplexer_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_2_io_inputs_1 = RegisterFile_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_2_io_inputs_0 = Multiplexer_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_3_io_configuration = Dispatch_3_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_3_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_3_io_inputs_3 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_3_io_inputs_2 = Multiplexer_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_3_io_inputs_1 = RegisterFile_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_3_io_inputs_0 = Multiplexer_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_4_io_configuration = Dispatch_3_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_4_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_4_io_inputs_3 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_4_io_inputs_2 = Multiplexer_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_4_io_inputs_1 = RegisterFile_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_4_io_inputs_0 = Multiplexer_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_5_io_configuration = Dispatch_3_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_5_io_inputs_1 = RegisterFile_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_5_io_inputs_0 = Multiplexer_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_6_io_configuration = Dispatch_3_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_6_io_inputs_1 = RegisterFile_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_6_io_inputs_0 = Multiplexer_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_7_io_configuration = Dispatch_3_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_7_io_inputs_1 = RegisterFile_26_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_7_io_inputs_0 = Multiplexer_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_configuration = Dispatch_4_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_8_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_8_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_configuration = Dispatch_4_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_9_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_9_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_configuration = Dispatch_4_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_10_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_10_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_configuration = Dispatch_4_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_11_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_11_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_configuration = Dispatch_4_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_12_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_12_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_configuration = Dispatch_4_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_13_io_inputs_5 = ConstUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_inputs_4 = Alu_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_inputs_3 = Multiplexer_25_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_inputs_2 = RegisterFile_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_13_io_inputs_0 = Multiplexer_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_14_io_configuration = Dispatch_4_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_14_io_inputs_1 = RegisterFile_29_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_14_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_15_io_configuration = Dispatch_4_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_15_io_inputs_1 = RegisterFile_30_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_15_io_inputs_0 = Multiplexer_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_16_io_configuration = Dispatch_4_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_16_io_inputs_1 = RegisterFile_31_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_16_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_17_io_configuration = Dispatch_4_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_17_io_inputs_1 = RegisterFile_32_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_17_io_inputs_0 = Multiplexer_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_configuration = Dispatch_5_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_18_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_18_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_configuration = Dispatch_5_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_19_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_19_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_configuration = Dispatch_5_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_20_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_20_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_configuration = Dispatch_5_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_21_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_21_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_configuration = Dispatch_5_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_22_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_22_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_configuration = Dispatch_5_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_23_io_inputs_5 = ConstUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_inputs_4 = Alu_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_inputs_3 = Multiplexer_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_inputs_2 = RegisterFile_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_23_io_inputs_0 = Multiplexer_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_24_io_configuration = Dispatch_5_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_24_io_inputs_1 = RegisterFile_35_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_24_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_25_io_configuration = Dispatch_5_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_25_io_inputs_1 = RegisterFile_36_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_25_io_inputs_0 = Multiplexer_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_26_io_configuration = Dispatch_5_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_26_io_inputs_1 = RegisterFile_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_26_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_27_io_configuration = Dispatch_5_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_27_io_inputs_1 = RegisterFile_38_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_27_io_inputs_0 = Multiplexer_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_configuration = Dispatch_6_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_28_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_28_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_configuration = Dispatch_6_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_29_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_29_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_configuration = Dispatch_6_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_30_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_30_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_configuration = Dispatch_6_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_31_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_31_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_configuration = Dispatch_6_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_32_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_32_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_configuration = Dispatch_6_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_33_io_inputs_5 = ConstUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_inputs_4 = Alu_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_inputs_3 = Multiplexer_45_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_inputs_2 = RegisterFile_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_33_io_inputs_0 = Multiplexer_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_34_io_configuration = Dispatch_6_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_34_io_inputs_1 = RegisterFile_41_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_34_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_35_io_configuration = Dispatch_6_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_35_io_inputs_1 = RegisterFile_42_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_35_io_inputs_0 = Multiplexer_29_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_36_io_configuration = Dispatch_6_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_36_io_inputs_1 = RegisterFile_43_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_36_io_inputs_0 = Multiplexer_30_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_37_io_configuration = Dispatch_6_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_37_io_inputs_1 = RegisterFile_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_37_io_inputs_0 = Multiplexer_31_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_configuration = Dispatch_7_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_38_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_38_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_configuration = Dispatch_7_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_39_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_39_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_configuration = Dispatch_7_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_40_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_40_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_configuration = Dispatch_7_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_41_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_41_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_configuration = Dispatch_7_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_42_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_42_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_configuration = Dispatch_7_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_43_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_inputs_4 = Alu_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_inputs_3 = Multiplexer_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_inputs_2 = RegisterFile_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_43_io_inputs_0 = Multiplexer_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_44_io_configuration = Dispatch_7_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_44_io_inputs_1 = RegisterFile_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_44_io_inputs_0 = Multiplexer_38_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_45_io_configuration = Dispatch_7_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_45_io_inputs_1 = RegisterFile_48_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_45_io_inputs_0 = Multiplexer_39_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_46_io_configuration = Dispatch_7_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_46_io_inputs_1 = RegisterFile_49_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_46_io_inputs_0 = Multiplexer_40_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_47_io_configuration = Dispatch_7_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_47_io_inputs_1 = RegisterFile_50_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_47_io_inputs_0 = Multiplexer_41_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_48_io_configuration = Dispatch_8_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_48_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_48_io_inputs_3 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_48_io_inputs_2 = RegisterFile_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_48_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_48_io_inputs_0 = Multiplexer_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_49_io_configuration = Dispatch_8_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_49_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_49_io_inputs_3 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_49_io_inputs_2 = RegisterFile_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_49_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_49_io_inputs_0 = Multiplexer_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_50_io_configuration = Dispatch_8_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_50_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_50_io_inputs_3 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_50_io_inputs_2 = RegisterFile_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_50_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_50_io_inputs_0 = Multiplexer_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_51_io_configuration = Dispatch_8_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_51_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_51_io_inputs_3 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_51_io_inputs_2 = RegisterFile_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_51_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_51_io_inputs_0 = Multiplexer_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_52_io_configuration = Dispatch_8_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_52_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_52_io_inputs_3 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_52_io_inputs_2 = RegisterFile_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_52_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_52_io_inputs_0 = Multiplexer_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_53_io_configuration = Dispatch_8_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_53_io_inputs_1 = RegisterFile_51_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_53_io_inputs_0 = Multiplexer_48_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_54_io_configuration = Dispatch_8_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_54_io_inputs_1 = RegisterFile_52_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_54_io_inputs_0 = Multiplexer_49_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_55_io_configuration = Dispatch_8_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_55_io_inputs_1 = RegisterFile_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_55_io_inputs_0 = Multiplexer_50_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_56_io_configuration = Dispatch_9_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_56_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_56_io_inputs_3 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_56_io_inputs_2 = Multiplexer_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_56_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_56_io_inputs_0 = Multiplexer_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_57_io_configuration = Dispatch_9_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_57_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_57_io_inputs_3 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_57_io_inputs_2 = Multiplexer_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_57_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_57_io_inputs_0 = Multiplexer_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_58_io_configuration = Dispatch_9_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_58_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_58_io_inputs_3 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_58_io_inputs_2 = Multiplexer_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_58_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_58_io_inputs_0 = Multiplexer_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_59_io_configuration = Dispatch_9_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_59_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_59_io_inputs_3 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_59_io_inputs_2 = Multiplexer_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_59_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_59_io_inputs_0 = Multiplexer_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_60_io_configuration = Dispatch_9_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_60_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_60_io_inputs_3 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_60_io_inputs_2 = Multiplexer_118_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_60_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_60_io_inputs_0 = Multiplexer_70_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_61_io_configuration = Dispatch_9_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_61_io_inputs_1 = RegisterFile_54_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_61_io_inputs_0 = Multiplexer_56_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_62_io_configuration = Dispatch_9_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_62_io_inputs_1 = RegisterFile_55_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_62_io_inputs_0 = Multiplexer_57_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_63_io_configuration = Dispatch_9_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_63_io_inputs_1 = RegisterFile_56_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_63_io_inputs_0 = Multiplexer_58_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_configuration = Dispatch_10_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_64_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_64_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_configuration = Dispatch_10_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_65_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_65_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_configuration = Dispatch_10_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_66_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_66_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_configuration = Dispatch_10_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_67_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_67_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_configuration = Dispatch_10_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_68_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_68_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_configuration = Dispatch_10_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_69_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_inputs_4 = Alu_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_inputs_3 = Multiplexer_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_inputs_2 = Multiplexer_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_inputs_1 = Multiplexer_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_69_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_70_io_configuration = Dispatch_10_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_70_io_inputs_1 = RegisterFile_59_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_70_io_inputs_0 = Multiplexer_64_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_71_io_configuration = Dispatch_10_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_71_io_inputs_1 = RegisterFile_60_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_71_io_inputs_0 = Multiplexer_65_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_72_io_configuration = Dispatch_10_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_72_io_inputs_1 = RegisterFile_61_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_72_io_inputs_0 = Multiplexer_66_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_73_io_configuration = Dispatch_10_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_73_io_inputs_1 = RegisterFile_62_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_73_io_inputs_0 = Multiplexer_67_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_configuration = Dispatch_11_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_74_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_74_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_configuration = Dispatch_11_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_75_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_75_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_configuration = Dispatch_11_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_76_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_76_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_configuration = Dispatch_11_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_77_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_77_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_configuration = Dispatch_11_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_78_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_78_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_configuration = Dispatch_11_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_79_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_inputs_4 = Alu_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_inputs_3 = Multiplexer_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_inputs_1 = Multiplexer_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_79_io_inputs_0 = Multiplexer_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_80_io_configuration = Dispatch_11_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_80_io_inputs_1 = RegisterFile_65_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_80_io_inputs_0 = Multiplexer_74_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_81_io_configuration = Dispatch_11_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_81_io_inputs_1 = RegisterFile_66_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_81_io_inputs_0 = Multiplexer_75_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_82_io_configuration = Dispatch_11_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_82_io_inputs_1 = RegisterFile_67_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_82_io_inputs_0 = Multiplexer_76_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_83_io_configuration = Dispatch_11_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_83_io_inputs_1 = RegisterFile_68_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_83_io_inputs_0 = Multiplexer_77_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_configuration = Dispatch_12_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_84_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_84_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_configuration = Dispatch_12_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_85_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_85_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_configuration = Dispatch_12_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_86_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_86_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_configuration = Dispatch_12_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_87_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_87_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_configuration = Dispatch_12_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_88_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_88_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_configuration = Dispatch_12_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_89_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_inputs_4 = Alu_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_inputs_3 = Multiplexer_148_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_inputs_2 = Multiplexer_34_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_inputs_1 = Multiplexer_100_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_89_io_inputs_0 = Multiplexer_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_90_io_configuration = Dispatch_12_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_90_io_inputs_1 = RegisterFile_71_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_90_io_inputs_0 = Multiplexer_84_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_91_io_configuration = Dispatch_12_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_91_io_inputs_1 = RegisterFile_72_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_91_io_inputs_0 = Multiplexer_85_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_92_io_configuration = Dispatch_12_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_92_io_inputs_1 = RegisterFile_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_92_io_inputs_0 = Multiplexer_86_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_93_io_configuration = Dispatch_12_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_93_io_inputs_1 = RegisterFile_74_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_93_io_inputs_0 = Multiplexer_87_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_configuration = Dispatch_13_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_94_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_94_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_configuration = Dispatch_13_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_95_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_95_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_configuration = Dispatch_13_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_96_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_96_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_configuration = Dispatch_13_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_97_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_97_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_configuration = Dispatch_13_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_98_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_98_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_configuration = Dispatch_13_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_99_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_inputs_4 = Alu_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_inputs_3 = Multiplexer_158_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_inputs_1 = Multiplexer_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_99_io_inputs_0 = Multiplexer_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_100_io_configuration = Dispatch_13_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_100_io_inputs_1 = RegisterFile_77_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_100_io_inputs_0 = Multiplexer_94_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_101_io_configuration = Dispatch_13_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_101_io_inputs_1 = RegisterFile_78_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_101_io_inputs_0 = Multiplexer_95_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_102_io_configuration = Dispatch_13_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_102_io_inputs_1 = RegisterFile_79_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_102_io_inputs_0 = Multiplexer_96_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_103_io_configuration = Dispatch_13_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_103_io_inputs_1 = RegisterFile_80_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_103_io_inputs_0 = Multiplexer_97_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_104_io_configuration = Dispatch_14_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_104_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_104_io_inputs_3 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_104_io_inputs_2 = Multiplexer_166_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_104_io_inputs_1 = Multiplexer_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_104_io_inputs_0 = Multiplexer_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_105_io_configuration = Dispatch_14_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_105_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_105_io_inputs_3 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_105_io_inputs_2 = Multiplexer_166_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_105_io_inputs_1 = Multiplexer_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_105_io_inputs_0 = Multiplexer_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_106_io_configuration = Dispatch_14_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_106_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_106_io_inputs_3 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_106_io_inputs_2 = Multiplexer_166_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_106_io_inputs_1 = Multiplexer_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_106_io_inputs_0 = Multiplexer_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_107_io_configuration = Dispatch_14_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_107_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_107_io_inputs_3 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_107_io_inputs_2 = Multiplexer_166_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_107_io_inputs_1 = Multiplexer_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_107_io_inputs_0 = Multiplexer_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_108_io_configuration = Dispatch_14_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_108_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_108_io_inputs_3 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_108_io_inputs_2 = Multiplexer_166_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_108_io_inputs_1 = Multiplexer_53_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_108_io_inputs_0 = Multiplexer_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_109_io_configuration = Dispatch_14_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_109_io_inputs_1 = RegisterFile_81_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_109_io_inputs_0 = Multiplexer_104_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_110_io_configuration = Dispatch_14_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_110_io_inputs_1 = RegisterFile_82_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_110_io_inputs_0 = Multiplexer_105_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_111_io_configuration = Dispatch_14_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_111_io_inputs_1 = RegisterFile_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_111_io_inputs_0 = Multiplexer_106_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_112_io_configuration = Dispatch_15_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_112_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_112_io_inputs_3 = LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_112_io_inputs_2 = Multiplexer_173_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_112_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_112_io_inputs_0 = Multiplexer_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_113_io_configuration = Dispatch_15_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_113_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_113_io_inputs_3 = LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_113_io_inputs_2 = Multiplexer_173_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_113_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_113_io_inputs_0 = Multiplexer_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_114_io_configuration = Dispatch_15_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_114_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_114_io_inputs_3 = LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_114_io_inputs_2 = Multiplexer_173_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_114_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_114_io_inputs_0 = Multiplexer_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_115_io_configuration = Dispatch_15_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_115_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_115_io_inputs_3 = LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_115_io_inputs_2 = Multiplexer_173_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_115_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_115_io_inputs_0 = Multiplexer_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_116_io_configuration = Dispatch_15_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_116_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_116_io_inputs_3 = LoadStoreUnit_4_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_116_io_inputs_2 = Multiplexer_173_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_116_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_116_io_inputs_0 = Multiplexer_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_117_io_configuration = Dispatch_15_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_117_io_inputs_1 = RegisterFile_84_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_117_io_inputs_0 = Multiplexer_112_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_118_io_configuration = Dispatch_15_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_118_io_inputs_1 = RegisterFile_85_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_118_io_inputs_0 = Multiplexer_113_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_119_io_configuration = Dispatch_15_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_119_io_inputs_1 = RegisterFile_86_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_119_io_inputs_0 = Multiplexer_114_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_configuration = Dispatch_16_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_120_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_120_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_configuration = Dispatch_16_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_121_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_121_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_configuration = Dispatch_16_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_122_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_122_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_configuration = Dispatch_16_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_123_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_123_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_configuration = Dispatch_16_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_124_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_124_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_configuration = Dispatch_16_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_125_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_inputs_4 = Alu_8_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_inputs_3 = Multiplexer_182_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_inputs_2 = Multiplexer_73_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_inputs_1 = Multiplexer_136_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_125_io_inputs_0 = Multiplexer_117_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_126_io_configuration = Dispatch_16_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_126_io_inputs_1 = RegisterFile_89_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_126_io_inputs_0 = Multiplexer_120_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_127_io_configuration = Dispatch_16_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_127_io_inputs_1 = RegisterFile_90_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_127_io_inputs_0 = Multiplexer_121_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_128_io_configuration = Dispatch_16_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_128_io_inputs_1 = RegisterFile_91_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_128_io_inputs_0 = Multiplexer_122_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_129_io_configuration = Dispatch_16_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_129_io_inputs_1 = RegisterFile_92_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_129_io_inputs_0 = Multiplexer_123_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_configuration = Dispatch_17_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_130_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_130_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_configuration = Dispatch_17_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_131_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_131_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_configuration = Dispatch_17_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_132_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_132_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_configuration = Dispatch_17_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_133_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_133_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_configuration = Dispatch_17_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_134_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_134_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_configuration = Dispatch_17_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_135_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_inputs_4 = Alu_9_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_inputs_3 = Multiplexer_192_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_inputs_2 = Multiplexer_83_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_inputs_1 = Multiplexer_146_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_135_io_inputs_0 = Multiplexer_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_136_io_configuration = Dispatch_17_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_136_io_inputs_1 = RegisterFile_95_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_136_io_inputs_0 = Multiplexer_130_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_137_io_configuration = Dispatch_17_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_137_io_inputs_1 = RegisterFile_96_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_137_io_inputs_0 = Multiplexer_131_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_138_io_configuration = Dispatch_17_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_138_io_inputs_1 = RegisterFile_97_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_138_io_inputs_0 = Multiplexer_132_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_139_io_configuration = Dispatch_17_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_139_io_inputs_1 = RegisterFile_98_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_139_io_inputs_0 = Multiplexer_133_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_configuration = Dispatch_18_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_140_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_140_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_configuration = Dispatch_18_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_141_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_141_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_configuration = Dispatch_18_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_142_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_142_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_configuration = Dispatch_18_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_143_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_143_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_configuration = Dispatch_18_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_144_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_144_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_configuration = Dispatch_18_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_145_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_inputs_4 = Alu_10_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_inputs_3 = Multiplexer_202_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_inputs_2 = Multiplexer_93_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_inputs_1 = Multiplexer_156_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_145_io_inputs_0 = Multiplexer_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_146_io_configuration = Dispatch_18_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_146_io_inputs_1 = RegisterFile_101_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_146_io_inputs_0 = Multiplexer_140_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_147_io_configuration = Dispatch_18_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_147_io_inputs_1 = RegisterFile_102_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_147_io_inputs_0 = Multiplexer_141_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_148_io_configuration = Dispatch_18_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_148_io_inputs_1 = RegisterFile_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_148_io_inputs_0 = Multiplexer_142_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_149_io_configuration = Dispatch_18_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_149_io_inputs_1 = RegisterFile_104_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_149_io_inputs_0 = Multiplexer_143_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_configuration = Dispatch_19_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_150_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_150_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_configuration = Dispatch_19_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_151_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_151_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_configuration = Dispatch_19_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_152_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_152_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_configuration = Dispatch_19_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_153_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_153_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_configuration = Dispatch_19_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_154_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_154_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_configuration = Dispatch_19_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_155_io_inputs_5 = ConstUnit_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_inputs_4 = Alu_11_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_inputs_3 = Multiplexer_212_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_inputs_2 = Multiplexer_103_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_inputs_1 = Multiplexer_165_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_155_io_inputs_0 = Multiplexer_147_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_156_io_configuration = Dispatch_19_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_156_io_inputs_1 = RegisterFile_107_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_156_io_inputs_0 = Multiplexer_150_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_157_io_configuration = Dispatch_19_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_157_io_inputs_1 = RegisterFile_108_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_157_io_inputs_0 = Multiplexer_151_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_158_io_configuration = Dispatch_19_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_158_io_inputs_1 = RegisterFile_109_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_158_io_inputs_0 = Multiplexer_152_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_159_io_configuration = Dispatch_19_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_159_io_inputs_1 = RegisterFile_110_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_159_io_inputs_0 = Multiplexer_153_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_160_io_configuration = Dispatch_20_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_160_io_inputs_4 = ConstUnit_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_160_io_inputs_3 = LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_160_io_inputs_2 = Multiplexer_221_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_160_io_inputs_1 = Multiplexer_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_160_io_inputs_0 = Multiplexer_157_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_161_io_configuration = Dispatch_20_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_161_io_inputs_4 = ConstUnit_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_161_io_inputs_3 = LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_161_io_inputs_2 = Multiplexer_221_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_161_io_inputs_1 = Multiplexer_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_161_io_inputs_0 = Multiplexer_157_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_162_io_configuration = Dispatch_20_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_162_io_inputs_4 = ConstUnit_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_162_io_inputs_3 = LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_162_io_inputs_2 = Multiplexer_221_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_162_io_inputs_1 = Multiplexer_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_162_io_inputs_0 = Multiplexer_157_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_163_io_configuration = Dispatch_20_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_163_io_inputs_4 = ConstUnit_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_163_io_inputs_3 = LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_163_io_inputs_2 = Multiplexer_221_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_163_io_inputs_1 = Multiplexer_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_163_io_inputs_0 = Multiplexer_157_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_164_io_configuration = Dispatch_20_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_164_io_inputs_4 = ConstUnit_17_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_164_io_inputs_3 = LoadStoreUnit_5_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_164_io_inputs_2 = Multiplexer_221_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_164_io_inputs_1 = Multiplexer_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_164_io_inputs_0 = Multiplexer_157_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_165_io_configuration = Dispatch_20_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_165_io_inputs_1 = RegisterFile_111_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_165_io_inputs_0 = Multiplexer_160_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_166_io_configuration = Dispatch_20_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_166_io_inputs_1 = RegisterFile_112_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_166_io_inputs_0 = Multiplexer_161_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_167_io_configuration = Dispatch_20_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_167_io_inputs_1 = RegisterFile_113_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_167_io_inputs_0 = Multiplexer_162_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_168_io_configuration = Dispatch_21_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_168_io_inputs_4 = ConstUnit_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_168_io_inputs_3 = LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_168_io_inputs_2 = Multiplexer_183_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_168_io_inputs_1 = Multiplexer_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_168_io_inputs_0 = RegisterFile_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_169_io_configuration = Dispatch_21_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_169_io_inputs_4 = ConstUnit_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_169_io_inputs_3 = LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_169_io_inputs_2 = Multiplexer_183_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_169_io_inputs_1 = Multiplexer_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_169_io_inputs_0 = RegisterFile_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_170_io_configuration = Dispatch_21_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_170_io_inputs_4 = ConstUnit_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_170_io_inputs_3 = LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_170_io_inputs_2 = Multiplexer_183_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_170_io_inputs_1 = Multiplexer_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_170_io_inputs_0 = RegisterFile_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_171_io_configuration = Dispatch_21_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_171_io_inputs_4 = ConstUnit_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_171_io_inputs_3 = LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_171_io_inputs_2 = Multiplexer_183_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_171_io_inputs_1 = Multiplexer_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_171_io_inputs_0 = RegisterFile_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_172_io_configuration = Dispatch_21_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_172_io_inputs_4 = ConstUnit_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_172_io_inputs_3 = LoadStoreUnit_6_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_172_io_inputs_2 = Multiplexer_183_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_172_io_inputs_1 = Multiplexer_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_172_io_inputs_0 = RegisterFile_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_173_io_configuration = Dispatch_21_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_173_io_inputs_1 = RegisterFile_114_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_173_io_inputs_0 = Multiplexer_168_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_174_io_configuration = Dispatch_21_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_174_io_inputs_1 = RegisterFile_115_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_174_io_inputs_0 = Multiplexer_169_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_175_io_configuration = Dispatch_21_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_175_io_inputs_1 = RegisterFile_116_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_175_io_inputs_0 = Multiplexer_170_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_configuration = Dispatch_22_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_176_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_176_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_configuration = Dispatch_22_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_177_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_177_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_configuration = Dispatch_22_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_178_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_178_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_configuration = Dispatch_22_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_179_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_179_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_configuration = Dispatch_22_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_180_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_180_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_configuration = Dispatch_22_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_181_io_inputs_5 = ConstUnit_19_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_inputs_4 = Alu_12_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_inputs_3 = Multiplexer_193_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_inputs_2 = Multiplexer_129_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_inputs_1 = RegisterFile_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_181_io_inputs_0 = Multiplexer_175_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_182_io_configuration = Dispatch_22_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_182_io_inputs_1 = RegisterFile_119_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_182_io_inputs_0 = Multiplexer_176_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_183_io_configuration = Dispatch_22_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_183_io_inputs_1 = RegisterFile_120_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_183_io_inputs_0 = Multiplexer_177_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_184_io_configuration = Dispatch_22_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_184_io_inputs_1 = RegisterFile_121_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_184_io_inputs_0 = Multiplexer_178_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_185_io_configuration = Dispatch_22_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_185_io_inputs_1 = RegisterFile_122_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_185_io_inputs_0 = Multiplexer_179_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_configuration = Dispatch_23_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_186_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_186_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_configuration = Dispatch_23_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_187_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_187_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_configuration = Dispatch_23_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_188_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_188_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_configuration = Dispatch_23_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_189_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_189_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_configuration = Dispatch_23_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_190_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_190_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_configuration = Dispatch_23_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_191_io_inputs_5 = ConstUnit_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_inputs_4 = Alu_13_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_inputs_3 = Multiplexer_203_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_inputs_2 = Multiplexer_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_inputs_1 = RegisterFile_16_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_191_io_inputs_0 = Multiplexer_185_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_192_io_configuration = Dispatch_23_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_192_io_inputs_1 = RegisterFile_125_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_192_io_inputs_0 = Multiplexer_186_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_193_io_configuration = Dispatch_23_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_193_io_inputs_1 = RegisterFile_126_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_193_io_inputs_0 = Multiplexer_187_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_194_io_configuration = Dispatch_23_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_194_io_inputs_1 = RegisterFile_127_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_194_io_inputs_0 = Multiplexer_188_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_195_io_configuration = Dispatch_23_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_195_io_inputs_1 = RegisterFile_128_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_195_io_inputs_0 = Multiplexer_189_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_configuration = Dispatch_24_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_196_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_196_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_configuration = Dispatch_24_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_197_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_197_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_configuration = Dispatch_24_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_198_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_198_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_configuration = Dispatch_24_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_199_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_199_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_configuration = Dispatch_24_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_200_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_200_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_configuration = Dispatch_24_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_201_io_inputs_5 = ConstUnit_21_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_inputs_4 = Alu_14_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_inputs_3 = Multiplexer_213_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_inputs_2 = Multiplexer_149_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_inputs_1 = RegisterFile_18_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_201_io_inputs_0 = Multiplexer_195_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_202_io_configuration = Dispatch_24_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_202_io_inputs_1 = RegisterFile_131_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_202_io_inputs_0 = Multiplexer_196_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_203_io_configuration = Dispatch_24_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_203_io_inputs_1 = RegisterFile_132_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_203_io_inputs_0 = Multiplexer_197_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_204_io_configuration = Dispatch_24_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_204_io_inputs_1 = RegisterFile_133_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_204_io_inputs_0 = Multiplexer_198_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_205_io_configuration = Dispatch_24_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_205_io_inputs_1 = RegisterFile_134_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_205_io_inputs_0 = Multiplexer_199_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_configuration = Dispatch_25_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_206_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_206_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_configuration = Dispatch_25_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_207_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_207_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_configuration = Dispatch_25_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_208_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_208_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_configuration = Dispatch_25_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_209_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_209_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_configuration = Dispatch_25_io_outs_11; // @[TopModule.scala 270:22]
  assign Multiplexer_210_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_210_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_configuration = Dispatch_25_io_outs_12; // @[TopModule.scala 270:22]
  assign Multiplexer_211_io_inputs_5 = ConstUnit_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_inputs_4 = Alu_15_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_inputs_3 = Multiplexer_222_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_inputs_2 = Multiplexer_159_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_inputs_1 = RegisterFile_20_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_211_io_inputs_0 = Multiplexer_205_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_212_io_configuration = Dispatch_25_io_outs_13; // @[TopModule.scala 270:22]
  assign Multiplexer_212_io_inputs_1 = RegisterFile_137_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_212_io_inputs_0 = Multiplexer_206_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_213_io_configuration = Dispatch_25_io_outs_14; // @[TopModule.scala 270:22]
  assign Multiplexer_213_io_inputs_1 = RegisterFile_138_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_213_io_inputs_0 = Multiplexer_207_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_214_io_configuration = Dispatch_25_io_outs_15; // @[TopModule.scala 270:22]
  assign Multiplexer_214_io_inputs_1 = RegisterFile_139_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_214_io_inputs_0 = Multiplexer_208_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_215_io_configuration = Dispatch_25_io_outs_16; // @[TopModule.scala 270:22]
  assign Multiplexer_215_io_inputs_1 = RegisterFile_140_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_215_io_inputs_0 = Multiplexer_209_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_216_io_configuration = Dispatch_26_io_outs_3; // @[TopModule.scala 270:22]
  assign Multiplexer_216_io_inputs_4 = ConstUnit_23_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_216_io_inputs_3 = LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_216_io_inputs_2 = Multiplexer_167_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_216_io_inputs_1 = RegisterFile_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_216_io_inputs_0 = Multiplexer_215_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_217_io_configuration = Dispatch_26_io_outs_4; // @[TopModule.scala 270:22]
  assign Multiplexer_217_io_inputs_4 = ConstUnit_23_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_217_io_inputs_3 = LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_217_io_inputs_2 = Multiplexer_167_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_217_io_inputs_1 = RegisterFile_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_217_io_inputs_0 = Multiplexer_215_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_218_io_configuration = Dispatch_26_io_outs_5; // @[TopModule.scala 270:22]
  assign Multiplexer_218_io_inputs_4 = ConstUnit_23_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_218_io_inputs_3 = LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_218_io_inputs_2 = Multiplexer_167_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_218_io_inputs_1 = RegisterFile_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_218_io_inputs_0 = Multiplexer_215_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_219_io_configuration = Dispatch_26_io_outs_6; // @[TopModule.scala 270:22]
  assign Multiplexer_219_io_inputs_4 = ConstUnit_23_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_219_io_inputs_3 = LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_219_io_inputs_2 = Multiplexer_167_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_219_io_inputs_1 = RegisterFile_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_219_io_inputs_0 = Multiplexer_215_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_220_io_configuration = Dispatch_26_io_outs_7; // @[TopModule.scala 270:22]
  assign Multiplexer_220_io_inputs_4 = ConstUnit_23_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_220_io_inputs_3 = LoadStoreUnit_7_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_220_io_inputs_2 = Multiplexer_167_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_220_io_inputs_1 = RegisterFile_22_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_220_io_inputs_0 = Multiplexer_215_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_221_io_configuration = Dispatch_26_io_outs_8; // @[TopModule.scala 270:22]
  assign Multiplexer_221_io_inputs_1 = RegisterFile_141_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_221_io_inputs_0 = Multiplexer_216_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_222_io_configuration = Dispatch_26_io_outs_9; // @[TopModule.scala 270:22]
  assign Multiplexer_222_io_inputs_1 = RegisterFile_142_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_222_io_inputs_0 = Multiplexer_217_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_223_io_configuration = Dispatch_26_io_outs_10; // @[TopModule.scala 270:22]
  assign Multiplexer_223_io_inputs_1 = RegisterFile_143_io_outs_0; // @[TopModule.scala 295:60]
  assign Multiplexer_223_io_inputs_0 = Multiplexer_218_io_outs_0; // @[TopModule.scala 295:60]
  assign ConstUnit_io_configuration = Dispatch_3_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_1_io_configuration = Dispatch_4_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_2_io_configuration = Dispatch_5_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_3_io_configuration = Dispatch_6_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_4_io_configuration = Dispatch_7_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_5_io_configuration = Dispatch_8_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_6_io_configuration = Dispatch_9_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_7_io_configuration = Dispatch_10_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_8_io_configuration = Dispatch_11_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_9_io_configuration = Dispatch_12_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_10_io_configuration = Dispatch_13_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_11_io_configuration = Dispatch_14_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_12_io_configuration = Dispatch_15_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_13_io_configuration = Dispatch_16_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_14_io_configuration = Dispatch_17_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_15_io_configuration = Dispatch_18_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_16_io_configuration = Dispatch_19_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_17_io_configuration = Dispatch_20_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_18_io_configuration = Dispatch_21_io_outs_11; // @[TopModule.scala 270:22]
  assign ConstUnit_19_io_configuration = Dispatch_22_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_20_io_configuration = Dispatch_23_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_21_io_configuration = Dispatch_24_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_22_io_configuration = Dispatch_25_io_outs_17; // @[TopModule.scala 270:22]
  assign ConstUnit_23_io_configuration = Dispatch_26_io_outs_11; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_clock = clock;
  assign LoadStoreUnit_reset = reset;
  assign LoadStoreUnit_io_configuration = Dispatch_3_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_io_en = MultiIIScheduleController_16_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_io_skewing = MultiIIScheduleController_16_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_io_streamIn_valid = io_streamInLSU_0_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_io_streamIn_bits = io_streamInLSU_0_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_io_len = io_lenLSU_0; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_io_streamOut_ready = io_streamOutLSU_0_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_io_base = io_baseLSU_0; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_io_start = io_startLSU_0; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_io_enqEn = io_enqEnLSU_0; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_io_deqEn = io_deqEnLSU_0; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_io_inputs_1 = Multiplexer_4_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_io_inputs_0 = Multiplexer_3_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_1_clock = clock;
  assign LoadStoreUnit_1_reset = reset;
  assign LoadStoreUnit_1_io_configuration = Dispatch_8_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_1_io_en = MultiIIScheduleController_17_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_1_io_skewing = MultiIIScheduleController_17_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_1_io_streamIn_valid = io_streamInLSU_1_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_1_io_streamIn_bits = io_streamInLSU_1_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_1_io_len = io_lenLSU_1; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_1_io_streamOut_ready = io_streamOutLSU_1_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_1_io_base = io_baseLSU_1; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_1_io_start = io_startLSU_1; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_1_io_enqEn = io_enqEnLSU_1; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_1_io_deqEn = io_deqEnLSU_1; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_1_io_inputs_1 = Multiplexer_52_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_1_io_inputs_0 = Multiplexer_51_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_2_clock = clock;
  assign LoadStoreUnit_2_reset = reset;
  assign LoadStoreUnit_2_io_configuration = Dispatch_9_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_2_io_en = MultiIIScheduleController_18_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_2_io_skewing = MultiIIScheduleController_18_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_2_io_streamIn_valid = io_streamInLSU_2_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_2_io_streamIn_bits = io_streamInLSU_2_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_2_io_len = io_lenLSU_2; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_2_io_streamOut_ready = io_streamOutLSU_2_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_2_io_base = io_baseLSU_2; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_2_io_start = io_startLSU_2; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_2_io_enqEn = io_enqEnLSU_2; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_2_io_deqEn = io_deqEnLSU_2; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_2_io_inputs_1 = Multiplexer_60_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_2_io_inputs_0 = Multiplexer_59_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_3_clock = clock;
  assign LoadStoreUnit_3_reset = reset;
  assign LoadStoreUnit_3_io_configuration = Dispatch_14_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_3_io_en = MultiIIScheduleController_19_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_3_io_skewing = MultiIIScheduleController_19_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_3_io_streamIn_valid = io_streamInLSU_3_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_3_io_streamIn_bits = io_streamInLSU_3_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_3_io_len = io_lenLSU_3; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_3_io_streamOut_ready = io_streamOutLSU_3_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_3_io_base = io_baseLSU_3; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_3_io_start = io_startLSU_3; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_3_io_enqEn = io_enqEnLSU_3; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_3_io_deqEn = io_deqEnLSU_3; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_3_io_inputs_1 = Multiplexer_108_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_3_io_inputs_0 = Multiplexer_107_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_4_clock = clock;
  assign LoadStoreUnit_4_reset = reset;
  assign LoadStoreUnit_4_io_configuration = Dispatch_15_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_4_io_en = MultiIIScheduleController_20_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_4_io_skewing = MultiIIScheduleController_20_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_4_io_streamIn_valid = io_streamInLSU_4_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_4_io_streamIn_bits = io_streamInLSU_4_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_4_io_len = io_lenLSU_4; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_4_io_streamOut_ready = io_streamOutLSU_4_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_4_io_base = io_baseLSU_4; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_4_io_start = io_startLSU_4; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_4_io_enqEn = io_enqEnLSU_4; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_4_io_deqEn = io_deqEnLSU_4; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_4_io_inputs_1 = Multiplexer_116_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_4_io_inputs_0 = Multiplexer_115_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_5_clock = clock;
  assign LoadStoreUnit_5_reset = reset;
  assign LoadStoreUnit_5_io_configuration = Dispatch_20_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_5_io_en = MultiIIScheduleController_21_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_5_io_skewing = MultiIIScheduleController_21_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_5_io_streamIn_valid = io_streamInLSU_5_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_5_io_streamIn_bits = io_streamInLSU_5_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_5_io_len = io_lenLSU_5; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_5_io_streamOut_ready = io_streamOutLSU_5_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_5_io_base = io_baseLSU_5; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_5_io_start = io_startLSU_5; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_5_io_enqEn = io_enqEnLSU_5; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_5_io_deqEn = io_deqEnLSU_5; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_5_io_inputs_1 = Multiplexer_164_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_5_io_inputs_0 = Multiplexer_163_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_6_clock = clock;
  assign LoadStoreUnit_6_reset = reset;
  assign LoadStoreUnit_6_io_configuration = Dispatch_21_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_6_io_en = MultiIIScheduleController_22_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_6_io_skewing = MultiIIScheduleController_22_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_6_io_streamIn_valid = io_streamInLSU_6_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_6_io_streamIn_bits = io_streamInLSU_6_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_6_io_len = io_lenLSU_6; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_6_io_streamOut_ready = io_streamOutLSU_6_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_6_io_base = io_baseLSU_6; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_6_io_start = io_startLSU_6; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_6_io_enqEn = io_enqEnLSU_6; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_6_io_deqEn = io_deqEnLSU_6; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_6_io_inputs_1 = Multiplexer_172_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_6_io_inputs_0 = Multiplexer_171_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_7_clock = clock;
  assign LoadStoreUnit_7_reset = reset;
  assign LoadStoreUnit_7_io_configuration = Dispatch_26_io_outs_12; // @[TopModule.scala 270:22]
  assign LoadStoreUnit_7_io_en = MultiIIScheduleController_23_io_valid; // @[TopModule.scala 210:17]
  assign LoadStoreUnit_7_io_skewing = MultiIIScheduleController_23_io_skewing; // @[TopModule.scala 211:22]
  assign LoadStoreUnit_7_io_streamIn_valid = io_streamInLSU_7_valid; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_7_io_streamIn_bits = io_streamInLSU_7_bits; // @[TopModule.scala 195:21]
  assign LoadStoreUnit_7_io_len = io_lenLSU_7; // @[TopModule.scala 190:16]
  assign LoadStoreUnit_7_io_streamOut_ready = io_streamOutLSU_7_ready; // @[TopModule.scala 196:22]
  assign LoadStoreUnit_7_io_base = io_baseLSU_7; // @[TopModule.scala 189:17]
  assign LoadStoreUnit_7_io_start = io_startLSU_7; // @[TopModule.scala 191:18]
  assign LoadStoreUnit_7_io_enqEn = io_enqEnLSU_7; // @[TopModule.scala 193:18]
  assign LoadStoreUnit_7_io_deqEn = io_deqEnLSU_7; // @[TopModule.scala 194:18]
  assign LoadStoreUnit_7_io_inputs_1 = Multiplexer_220_io_outs_0; // @[TopModule.scala 295:60]
  assign LoadStoreUnit_7_io_inputs_0 = Multiplexer_219_io_outs_0[5:0]; // @[TopModule.scala 295:60]
  assign MultiIIScheduleController_16_clock = clock;
  assign MultiIIScheduleController_16_reset = reset;
  assign MultiIIScheduleController_16_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_16_io_schedules_0 = Dispatch_io_outs_128; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_1 = Dispatch_io_outs_129; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_2 = Dispatch_io_outs_130; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_3 = Dispatch_io_outs_131; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_4 = Dispatch_io_outs_132; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_5 = Dispatch_io_outs_133; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_6 = Dispatch_io_outs_134; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_schedules_7 = Dispatch_io_outs_135; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_16_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_17_clock = clock;
  assign MultiIIScheduleController_17_reset = reset;
  assign MultiIIScheduleController_17_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_17_io_schedules_0 = Dispatch_io_outs_136; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_1 = Dispatch_io_outs_137; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_2 = Dispatch_io_outs_138; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_3 = Dispatch_io_outs_139; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_4 = Dispatch_io_outs_140; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_5 = Dispatch_io_outs_141; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_6 = Dispatch_io_outs_142; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_schedules_7 = Dispatch_io_outs_143; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_17_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_18_clock = clock;
  assign MultiIIScheduleController_18_reset = reset;
  assign MultiIIScheduleController_18_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_18_io_schedules_0 = Dispatch_io_outs_144; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_1 = Dispatch_io_outs_145; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_2 = Dispatch_io_outs_146; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_3 = Dispatch_io_outs_147; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_4 = Dispatch_io_outs_148; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_5 = Dispatch_io_outs_149; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_6 = Dispatch_io_outs_150; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_schedules_7 = Dispatch_io_outs_151; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_18_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_19_clock = clock;
  assign MultiIIScheduleController_19_reset = reset;
  assign MultiIIScheduleController_19_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_19_io_schedules_0 = Dispatch_io_outs_152; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_1 = Dispatch_io_outs_153; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_2 = Dispatch_io_outs_154; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_3 = Dispatch_io_outs_155; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_4 = Dispatch_io_outs_156; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_5 = Dispatch_io_outs_157; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_6 = Dispatch_io_outs_158; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_schedules_7 = Dispatch_io_outs_159; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_19_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_20_clock = clock;
  assign MultiIIScheduleController_20_reset = reset;
  assign MultiIIScheduleController_20_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_20_io_schedules_0 = Dispatch_io_outs_160; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_1 = Dispatch_io_outs_161; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_2 = Dispatch_io_outs_162; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_3 = Dispatch_io_outs_163; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_4 = Dispatch_io_outs_164; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_5 = Dispatch_io_outs_165; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_6 = Dispatch_io_outs_166; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_schedules_7 = Dispatch_io_outs_167; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_20_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_21_clock = clock;
  assign MultiIIScheduleController_21_reset = reset;
  assign MultiIIScheduleController_21_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_21_io_schedules_0 = Dispatch_io_outs_168; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_1 = Dispatch_io_outs_169; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_2 = Dispatch_io_outs_170; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_3 = Dispatch_io_outs_171; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_4 = Dispatch_io_outs_172; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_5 = Dispatch_io_outs_173; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_6 = Dispatch_io_outs_174; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_schedules_7 = Dispatch_io_outs_175; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_21_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_22_clock = clock;
  assign MultiIIScheduleController_22_reset = reset;
  assign MultiIIScheduleController_22_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_22_io_schedules_0 = Dispatch_io_outs_176; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_1 = Dispatch_io_outs_177; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_2 = Dispatch_io_outs_178; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_3 = Dispatch_io_outs_179; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_4 = Dispatch_io_outs_180; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_5 = Dispatch_io_outs_181; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_6 = Dispatch_io_outs_182; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_schedules_7 = Dispatch_io_outs_183; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_22_io_II = io_II; // @[TopModule.scala 206:38]
  assign MultiIIScheduleController_23_clock = clock;
  assign MultiIIScheduleController_23_reset = reset;
  assign MultiIIScheduleController_23_io_en = io_en; // @[TopModule.scala 205:38]
  assign MultiIIScheduleController_23_io_schedules_0 = Dispatch_io_outs_184; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_1 = Dispatch_io_outs_185; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_2 = Dispatch_io_outs_186; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_3 = Dispatch_io_outs_187; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_4 = Dispatch_io_outs_188; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_5 = Dispatch_io_outs_189; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_6 = Dispatch_io_outs_190; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_schedules_7 = Dispatch_io_outs_191; // @[TopModule.scala 208:50]
  assign MultiIIScheduleController_23_io_II = io_II; // @[TopModule.scala 206:38]
  assign configControllers_0_clock = clock;
  assign configControllers_0_reset = reset;
  assign configControllers_0_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_0_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_0_io_inConfig = topDispatch_io_outs_0; // @[TopModule.scala 280:38]
  assign Dispatch_1_io_configuration = configControllers_0_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_1_clock = clock;
  assign configControllers_1_reset = reset;
  assign configControllers_1_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_1_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_1_io_inConfig = topDispatch_io_outs_1; // @[TopModule.scala 280:38]
  assign Dispatch_2_io_configuration = configControllers_1_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_2_clock = clock;
  assign configControllers_2_reset = reset;
  assign configControllers_2_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_2_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_2_io_inConfig = topDispatch_io_outs_2; // @[TopModule.scala 280:38]
  assign Dispatch_3_io_configuration = configControllers_2_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_3_clock = clock;
  assign configControllers_3_reset = reset;
  assign configControllers_3_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_3_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_3_io_inConfig = topDispatch_io_outs_3; // @[TopModule.scala 280:38]
  assign Dispatch_4_io_configuration = configControllers_3_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_4_clock = clock;
  assign configControllers_4_reset = reset;
  assign configControllers_4_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_4_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_4_io_inConfig = topDispatch_io_outs_4; // @[TopModule.scala 280:38]
  assign Dispatch_5_io_configuration = configControllers_4_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_5_clock = clock;
  assign configControllers_5_reset = reset;
  assign configControllers_5_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_5_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_5_io_inConfig = topDispatch_io_outs_5; // @[TopModule.scala 280:38]
  assign Dispatch_6_io_configuration = configControllers_5_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_6_clock = clock;
  assign configControllers_6_reset = reset;
  assign configControllers_6_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_6_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_6_io_inConfig = topDispatch_io_outs_6; // @[TopModule.scala 280:38]
  assign Dispatch_7_io_configuration = configControllers_6_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_7_clock = clock;
  assign configControllers_7_reset = reset;
  assign configControllers_7_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_7_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_7_io_inConfig = topDispatch_io_outs_7; // @[TopModule.scala 280:38]
  assign Dispatch_8_io_configuration = configControllers_7_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_8_clock = clock;
  assign configControllers_8_reset = reset;
  assign configControllers_8_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_8_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_8_io_inConfig = topDispatch_io_outs_8; // @[TopModule.scala 280:38]
  assign Dispatch_9_io_configuration = configControllers_8_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_9_clock = clock;
  assign configControllers_9_reset = reset;
  assign configControllers_9_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_9_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_9_io_inConfig = topDispatch_io_outs_9; // @[TopModule.scala 280:38]
  assign Dispatch_10_io_configuration = configControllers_9_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_10_clock = clock;
  assign configControllers_10_reset = reset;
  assign configControllers_10_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_10_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_10_io_inConfig = topDispatch_io_outs_10; // @[TopModule.scala 280:38]
  assign Dispatch_11_io_configuration = configControllers_10_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_11_clock = clock;
  assign configControllers_11_reset = reset;
  assign configControllers_11_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_11_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_11_io_inConfig = topDispatch_io_outs_11; // @[TopModule.scala 280:38]
  assign Dispatch_12_io_configuration = configControllers_11_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_12_clock = clock;
  assign configControllers_12_reset = reset;
  assign configControllers_12_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_12_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_12_io_inConfig = topDispatch_io_outs_12; // @[TopModule.scala 280:38]
  assign Dispatch_13_io_configuration = configControllers_12_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_13_clock = clock;
  assign configControllers_13_reset = reset;
  assign configControllers_13_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_13_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_13_io_inConfig = topDispatch_io_outs_13; // @[TopModule.scala 280:38]
  assign Dispatch_14_io_configuration = configControllers_13_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_14_clock = clock;
  assign configControllers_14_reset = reset;
  assign configControllers_14_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_14_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_14_io_inConfig = topDispatch_io_outs_14; // @[TopModule.scala 280:38]
  assign Dispatch_15_io_configuration = configControllers_14_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_15_clock = clock;
  assign configControllers_15_reset = reset;
  assign configControllers_15_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_15_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_15_io_inConfig = topDispatch_io_outs_15; // @[TopModule.scala 280:38]
  assign Dispatch_16_io_configuration = configControllers_15_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_16_clock = clock;
  assign configControllers_16_reset = reset;
  assign configControllers_16_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_16_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_16_io_inConfig = topDispatch_io_outs_16; // @[TopModule.scala 280:38]
  assign Dispatch_17_io_configuration = configControllers_16_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_17_clock = clock;
  assign configControllers_17_reset = reset;
  assign configControllers_17_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_17_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_17_io_inConfig = topDispatch_io_outs_17; // @[TopModule.scala 280:38]
  assign Dispatch_18_io_configuration = configControllers_17_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_18_clock = clock;
  assign configControllers_18_reset = reset;
  assign configControllers_18_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_18_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_18_io_inConfig = topDispatch_io_outs_18; // @[TopModule.scala 280:38]
  assign Dispatch_19_io_configuration = configControllers_18_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_19_clock = clock;
  assign configControllers_19_reset = reset;
  assign configControllers_19_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_19_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_19_io_inConfig = topDispatch_io_outs_19; // @[TopModule.scala 280:38]
  assign Dispatch_20_io_configuration = configControllers_19_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_20_clock = clock;
  assign configControllers_20_reset = reset;
  assign configControllers_20_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_20_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_20_io_inConfig = topDispatch_io_outs_20; // @[TopModule.scala 280:38]
  assign Dispatch_21_io_configuration = configControllers_20_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_21_clock = clock;
  assign configControllers_21_reset = reset;
  assign configControllers_21_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_21_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_21_io_inConfig = topDispatch_io_outs_21; // @[TopModule.scala 280:38]
  assign Dispatch_22_io_configuration = configControllers_21_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_22_clock = clock;
  assign configControllers_22_reset = reset;
  assign configControllers_22_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_22_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_22_io_inConfig = topDispatch_io_outs_22; // @[TopModule.scala 280:38]
  assign Dispatch_23_io_configuration = configControllers_22_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_23_clock = clock;
  assign configControllers_23_reset = reset;
  assign configControllers_23_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_23_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_23_io_inConfig = topDispatch_io_outs_23; // @[TopModule.scala 280:38]
  assign Dispatch_24_io_configuration = configControllers_23_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_24_clock = clock;
  assign configControllers_24_reset = reset;
  assign configControllers_24_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_24_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_24_io_inConfig = topDispatch_io_outs_24; // @[TopModule.scala 280:38]
  assign Dispatch_25_io_configuration = configControllers_24_io_outConfig; // @[TopModule.scala 273:31]
  assign configControllers_25_clock = clock;
  assign configControllers_25_reset = reset;
  assign configControllers_25_io_en = io_enConfig; // @[TopModule.scala 264:28]
  assign configControllers_25_io_II = io_II; // @[TopModule.scala 263:28]
  assign configControllers_25_io_inConfig = topDispatch_io_outs_25; // @[TopModule.scala 280:38]
  assign Dispatch_26_io_configuration = configControllers_25_io_outConfig; // @[TopModule.scala 273:31]
  assign topDispatch_io_configuration = io_configuration; // @[TopModule.scala 278:32]
endmodule
